* SPICE3 file created from total.ext - technology: sky130A
VVSS VSS 0 0
VVCC VCC VSS 3.3

VINP INP INN sin(0 shift 4e6)
VINN INN VSS VMEAN

x1 VCC VSS INP INN VOUT total

**** begin user architecture code

.option chgtol=4e-16 method=gear

.param VMEAN = 0
.param shift = 2m

**** interactive sim
.control
run
save all
tran 20n 2u
plot ((inp-inn)*100)+1.65 vout 
.endc


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/ff.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/ff/specialized_cells.spice


.subckt total VCC VSS INP INN VOUT
X0 m1_6795_368# diff_to_single_ended_1/v VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.143 ps=1.06 w=0.5 l=0.5
X1 VSS current_source_0/li_1035_74# VSS sky130_fd_pr__res_generic_nd__hv w=0.415 l=5.8
X2 current_source_0/li_1035_74# VSS VSS sky130_fd_pr__res_generic_nd__hv w=0.415 l=5.8
X3 folded_cascode_0/Vb3 current_source_0/li_1085_2889# current_source_0/m1_737_3994# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.5 w=3 l=2
X4 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=2
X5 current_source_0/li_226_2694# current_source_0/li_1085_2889# current_source_0/m1_1325_3826# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.5 w=3 l=2
X6 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=2
X7 current_source_0/m1_737_3994# current_source_0/li_1085_2889# folded_cascode_0/Vb3 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.5 as=0.87 ps=6.58 w=3 l=2
X8 current_source_0/m1_1325_3826# current_source_0/li_1085_2889# current_source_0/li_226_2694# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.5 as=0.87 ps=6.58 w=3 l=2
X9 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=2
X10 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.856 pd=6.36 as=0.856 ps=6.36 w=3 l=2
X11 VCC current_source_0/a_798_3689# current_source_0/m1_737_3994# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=1.16 ps=8.66 w=4 l=2
X12 input_stage_0/Vb5 folded_cascode_0/Vb3 folded_cascode_0/Vb3 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.39 as=0.58 ps=4.58 w=2 l=0.5
X13 VCC current_source_0/a_798_3689# current_source_0/m1_1325_3826# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=1.16 ps=8.66 w=4 l=2
X14 VCC current_source_0/a_798_3689# current_source_0/a_798_3689# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.911 ps=6.78 w=4 l=2
X15 current_source_0/a_798_3689# current_source_0/a_798_3689# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.911 pd=6.78 as=0.998 ps=7.37 w=4 l=2
X16 current_source_0/m1_1913_2070# current_source_0/li_805_1641# current_source_0/li_1035_74# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.55 pd=11.2 as=2.49 ps=18.4 w=8 l=2
X17 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.28 pd=17 as=2.28 ps=17 w=8 l=2
X18 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.28 pd=17 as=2.28 ps=17 w=8 l=2
X19 current_source_0/li_1035_74# current_source_0/li_805_1641# current_source_0/m1_1913_2070# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.49 pd=18.4 as=1.55 ps=11.2 w=8 l=2
X20 current_source_0/li_1085_2889# current_source_0/li_1085_2889# current_source_0/a_798_3689# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.684 ps=5.09 w=3 l=2
X21 current_source_0/a_798_3689# current_source_0/li_1085_2889# current_source_0/li_1085_2889# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.684 pd=5.09 as=0.87 ps=6.58 w=3 l=2
X22 folded_cascode_0/Vb2 current_source_0/li_226_2694# current_source_0/m1_737_1534# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X23 current_source_0/li_226_2694# current_source_0/li_226_2694# current_source_0/li_805_1641# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X24 current_source_0/li_1085_2889# current_source_0/li_226_2694# current_source_0/m1_1913_2070# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.773 ps=5.62 w=4 l=2
X25 input_stage_0/Vb5 input_stage_0/Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.77 as=1.14 ps=8.49 w=4 l=0.5
X26 current_source_0/m1_1913_2070# current_source_0/li_226_2694# current_source_0/li_1085_2889# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.773 pd=5.62 as=0.58 ps=4.29 w=4 l=2
X27 current_source_0/m1_1325_3826# current_source_0/a_798_3689# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.66 as=0.998 ps=7.37 w=4 l=2
X28 current_source_0/li_805_1641# current_source_0/li_226_2694# current_source_0/li_226_2694# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X29 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.14 ps=8.49 w=4 l=2
X30 current_source_0/m1_737_3994# current_source_0/a_798_3689# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.66 as=0.998 ps=7.37 w=4 l=2
X31 current_source_0/li_805_1641# current_source_0/li_805_1641# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.14 ps=8.49 w=4 l=2
X32 VSS current_source_0/li_805_1641# current_source_0/li_805_1641# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.16 ps=8.58 w=4 l=2
X33 VSS current_source_0/li_805_1641# current_source_0/m1_737_1534# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.16 ps=8.58 w=4 l=2
X34 current_source_0/m1_737_1534# current_source_0/li_805_1641# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.14 ps=8.49 w=4 l=2
X35 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.14 ps=8.49 w=4 l=2
X36 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=3.77 pd=28 as=3.77 ps=28 w=13.2 l=0.5
X37 current_source_0/m1_737_1534# current_source_0/li_226_2694# folded_cascode_0/Vb2 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X38 VSS current_source_0/m1_151_2991# current_source_0/a_798_3689# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.16 ps=8.58 w=4 l=2
X39 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=3.77 pd=28 as=3.77 ps=28 w=13.2 l=0.5
X40 VSS current_source_0/li_226_2694# current_source_0/m1_151_2991# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.16 ps=8.58 w=4 l=2
X41 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=3.77 pd=28 as=3.77 ps=28 w=13.2 l=0.5
X42 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.748 pd=5.53 as=0.748 ps=5.53 w=3 l=2
X43 VCC cmfb_block_0/Vb1 cmfb_block_0/Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2 pd=14.7 as=2.32 ps=16.6 w=8 l=0.5
X44 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.54 pd=11.5 as=1.54 ps=11.5 w=5.4 l=0.5
X45 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2 pd=14.7 as=2 ps=14.7 w=8 l=0.5
X46 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.748 pd=5.53 as=0.748 ps=5.53 w=3 l=2
X47 cmfb_block_0/Vb1 folded_cascode_0/Vb2 folded_cascode_0/Vb2 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=0.5
X48 VSS current_source_0/li_1035_74# VSS sky130_fd_pr__res_generic_nd__hv w=0.415 l=5.8
X49 VCC current_source_0/li_226_2694# current_source_0/m1_151_2991# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.748 pd=5.53 as=0.87 ps=6.58 w=3 l=2
X50 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2 pd=14.7 as=2 ps=14.7 w=8 l=0.5
X51 current_source_0/li_1035_74# VSS VSS sky130_fd_pr__res_generic_nd__hv w=0.415 l=5.8
X52 cmfb_block_0/m1_3052_n816# cmfb_block_0/VREF cmfb_block_0/CMFB VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.887 pd=6.8 as=1.16 ps=8.58 w=4 l=0.5
X53 cmfb_block_0/CMFB cmfb_block_0/VREF cmfb_block_0/m1_3052_n816# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.887 ps=6.8 w=4 l=0.5
X54 cmfb_block_0/a_2761_n1936# cmfb_block_0/IN cmfb_block_0/m1_3637_198# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.887 ps=6.8 w=4 l=0.5
X55 VCC cmfb_block_0/Vb1 cmfb_block_0/m1_3637_198# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.111 ps=0.85 w=0.5 l=0.5
X56 cmfb_block_0/m1_3052_n816# cmfb_block_0/Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=0.85 as=0.125 ps=0.922 w=0.5 l=0.5
X57 cmfb_block_0/m1_3637_198# cmfb_block_0/IN cmfb_block_0/a_2761_n1936# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.887 pd=6.8 as=1.16 ps=8.58 w=4 l=0.5
X58 VCC cmfb_block_0/Vb1 cmfb_block_0/m1_3052_n816# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.111 ps=0.85 w=0.5 l=0.5
X59 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.125 ps=0.922 w=0.5 l=1.5
X60 cmfb_block_0/m1_3637_198# cmfb_block_0/VREF cmfb_block_0/CMFB VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.887 pd=6.8 as=1.16 ps=8.58 w=4 l=0.5
X61 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.125 ps=0.922 w=0.5 l=1.5
X62 cmfb_block_0/m1_3637_198# cmfb_block_0/Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=0.85 as=0.125 ps=0.922 w=0.5 l=0.5
X63 cmfb_block_0/CMFB cmfb_block_0/VREF cmfb_block_0/m1_3637_198# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.887 ps=6.8 w=4 l=0.5
X64 cmfb_block_0/a_2761_n1936# cmfb_block_0/IP cmfb_block_0/m1_3052_n816# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.887 ps=6.8 w=4 l=0.5
X65 cmfb_block_0/m1_3052_n816# cmfb_block_0/IP cmfb_block_0/a_2761_n1936# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.887 pd=6.8 as=1.16 ps=8.58 w=4 l=0.5
X66 VSS cmfb_block_0/CMFB cmfb_block_0/CMFB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.145 ps=1.58 w=0.5 l=1
X67 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.143 ps=1.06 w=0.5 l=0.5
X68 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.143 ps=1.06 w=0.5 l=0.5
X69 VSS cmfb_block_0/a_2761_n1936# cmfb_block_0/a_2761_n1936# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.145 ps=1.58 w=0.5 l=1
X70 cmfb_block_0/CMFB cmfb_block_0/CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.143 ps=1.06 w=0.5 l=1
X71 cmfb_block_0/a_2761_n1936# cmfb_block_0/a_2761_n1936# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.143 ps=1.06 w=0.5 l=1
X72 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=1.5
X73 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=1.5
X74 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=1.5
X75 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=1.5
X76 cmfb_block_0/CMFB VSS sky130_fd_pr__cap_mim_m3_1 l=6 w=7.1
X77 VOUT m1_6795_368# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=2.49 ps=18.4 w=10 l=0.5
X78 m1_6795_368# diff_to_single_ended_1/v VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.25 ps=9.22 w=5 l=0.5
X79 diff_to_single_ended_1/a_n296_n44# cmfb_block_0/IN diff_to_single_ended_1/li_n130_n833# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.464 ps=4.01 w=2 l=0.5
X80 VSS input_stage_0/Vb5 diff_to_single_ended_1/li_n130_n833# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.116 ps=1 w=0.5 l=0.5
X81 diff_to_single_ended_1/li_n130_n833# input_stage_0/Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.116 pd=1 as=0.143 ps=1.06 w=0.5 l=0.5
X82 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.143 ps=1.06 w=0.5 l=2
X83 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.143 ps=1.06 w=0.5 l=2
X84 diff_to_single_ended_1/li_n130_n833# input_stage_0/Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.116 pd=1 as=0.143 ps=1.06 w=0.5 l=0.5
X85 VSS input_stage_0/Vb5 diff_to_single_ended_1/li_n130_n833# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.116 ps=1 w=0.5 l=0.5
X86 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.571 pd=4.24 as=0.571 ps=4.24 w=2 l=2
X87 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.571 pd=4.24 as=0.571 ps=4.24 w=2 l=2
X88 VCC diff_to_single_ended_1/a_n296_n44# diff_to_single_ended_1/a_n296_n44# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.145 ps=1.58 w=0.5 l=1
X89 diff_to_single_ended_1/v diff_to_single_ended_1/a_n296_n44# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.125 ps=0.922 w=0.5 l=1
X90 VCC diff_to_single_ended_1/a_n296_n44# diff_to_single_ended_1/v VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.145 ps=1.58 w=0.5 l=1
X91 diff_to_single_ended_1/a_n296_n44# diff_to_single_ended_1/a_n296_n44# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.125 ps=0.922 w=0.5 l=1
X92 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.125 ps=0.922 w=0.5 l=0.5
X93 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.125 pd=0.922 as=0.125 ps=0.922 w=0.5 l=0.5
X94 diff_to_single_ended_1/li_n130_n833# cmfb_block_0/IP diff_to_single_ended_1/v VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=4.01 as=0.58 ps=4.58 w=2 l=0.5
X95 diff_to_single_ended_1/v cmfb_block_0/IP diff_to_single_ended_1/li_n130_n833# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.464 ps=4.01 w=2 l=0.5
X96 diff_to_single_ended_1/li_n130_n833# cmfb_block_0/IN diff_to_single_ended_1/a_n296_n44# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=4.01 as=0.58 ps=4.58 w=2 l=0.5
X97 cmfb_block_0/VREF VCC VCC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=9.03 as=19.4 ps=163 w=4 l=0.5
X98 input_stage_0/N2 cmfb_block_0/Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.93 as=0.998 ps=7.37 w=4 l=0.5
X99 VCC cmfb_block_0/Vb1 input_stage_0/N2 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=1.16 ps=8.93 w=4 l=0.5
X100 input_stage_0/N3 folded_cascode_0/Vb3 cmfb_block_0/IP VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.39 as=0.58 ps=4.58 w=2 l=0.5
X101 input_stage_0/N3 cmfb_block_0/CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.77 as=1.14 ps=8.49 w=4 l=0.5
X102 VCC cmfb_block_0/Vb1 input_stage_0/N1 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=1.16 ps=8.93 w=4 l=0.5
X103 input_stage_0/N4 cmfb_block_0/CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.77 as=1.14 ps=8.49 w=4 l=0.5
X104 VSS cmfb_block_0/CMFB input_stage_0/N4 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.16 ps=8.77 w=4 l=0.5
X105 VSS cmfb_block_0/CMFB input_stage_0/N3 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.16 ps=8.77 w=4 l=0.5
X106 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.14 ps=8.49 w=4 l=0.5
X107 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.14 pd=8.49 as=1.14 ps=8.49 w=4 l=0.5
X108 cmfb_block_0/IN folded_cascode_0/Vb2 input_stage_0/N2 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.23 w=1 l=0.5
X109 input_stage_0/N2 folded_cascode_0/Vb2 cmfb_block_0/IN VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.23 as=0.145 ps=1.29 w=1 l=0.5
X110 input_stage_0/N1 folded_cascode_0/Vb2 cmfb_block_0/IP VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.23 as=0.29 ps=2.58 w=1 l=0.5
X111 cmfb_block_0/IP folded_cascode_0/Vb2 input_stage_0/N1 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.23 w=1 l=0.5
X112 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.571 pd=4.24 as=0.571 ps=4.24 w=2 l=0.5
X113 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.571 pd=4.24 as=0.571 ps=4.24 w=2 l=0.5
X114 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.249 pd=1.84 as=0.249 ps=1.84 w=1 l=0.5
X115 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.249 pd=1.84 as=0.249 ps=1.84 w=1 l=0.5
X116 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=0.5
X117 input_stage_0/N4 folded_cascode_0/Vb3 cmfb_block_0/IN VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.39 as=0.29 ps=2.29 w=2 l=0.5
X118 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.998 pd=7.37 as=0.998 ps=7.37 w=4 l=0.5
X119 cmfb_block_0/IP folded_cascode_0/Vb3 input_stage_0/N3 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.39 w=2 l=0.5
X120 cmfb_block_0/IN folded_cascode_0/Vb3 input_stage_0/N4 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.39 w=2 l=0.5
X121 input_stage_0/N1 cmfb_block_0/Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.93 as=0.998 ps=7.37 w=4 l=0.5
X122 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2 pd=14.7 as=2 ps=14.7 w=8 l=0.5
X123 input_stage_0/m1_n402_n3947# input_stage_0/Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=0.824 as=0.143 ps=1.06 w=0.5 l=0.5
X124 input_stage_0/m1_n402_n3947# input_stage_0/Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=0.824 as=0.143 ps=1.06 w=0.5 l=0.5
X125 VSS input_stage_0/Vb5 input_stage_0/m1_n402_n3947# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.111 ps=0.824 w=0.5 l=0.5
X126 VSS input_stage_0/Vb5 input_stage_0/m1_n402_n3947# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.111 ps=0.824 w=0.5 l=0.5
X127 input_stage_0/N4 INN input_stage_0/m1_n402_90# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.8 ps=13.3 w=8 l=0.5
X128 input_stage_0/N3 INP input_stage_0/m1_n402_90# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.8 ps=13.3 w=8 l=0.5
X129 input_stage_0/m1_n402_90# INN input_stage_0/N4 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.8 pd=13.3 as=2.32 ps=16.6 w=8 l=0.5
X130 input_stage_0/m1_n402_90# INP input_stage_0/N3 VCC sky130_fd_pr__pfet_g5v0d10v5 ad=1.8 pd=13.3 as=2.32 ps=16.6 w=8 l=0.5
X131 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.28 pd=17 as=2.28 ps=17 w=8 l=0.5
X132 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.143 ps=1.06 w=0.5 l=0.5
X133 input_stage_0/m1_n402_90# cmfb_block_0/Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.226 pd=1.67 as=0.249 ps=1.84 w=1 l=0.5
X134 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.28 pd=17 as=2.28 ps=17 w=8 l=0.5
X135 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.143 pd=1.06 as=0.143 ps=1.06 w=0.5 l=0.5
X136 input_stage_0/m1_n402_90# cmfb_block_0/Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.226 pd=1.67 as=0.249 ps=1.84 w=1 l=0.5
X137 VCC cmfb_block_0/Vb1 input_stage_0/m1_n402_90# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.249 pd=1.84 as=0.226 ps=1.67 w=1 l=0.5
X138 VCC cmfb_block_0/Vb1 input_stage_0/m1_n402_90# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.249 pd=1.84 as=0.226 ps=1.67 w=1 l=0.5
X139 input_stage_0/m1_n402_n3947# INN input_stage_0/N2 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.77 pd=13.2 as=2.32 ps=16.6 w=8 l=0.5
X140 input_stage_0/N2 INN input_stage_0/m1_n402_n3947# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.77 ps=13.2 w=8 l=0.5
X141 input_stage_0/m1_n402_n3947# INP input_stage_0/N1 VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.77 pd=13.2 as=2.32 ps=16.6 w=8 l=0.5
X142 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.249 pd=1.84 as=0.249 ps=1.84 w=1 l=0.5
X143 input_stage_0/N1 INP input_stage_0/m1_n402_n3947# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.77 ps=13.2 w=8 l=0.5
X144 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.249 pd=1.84 as=0.249 ps=1.84 w=1 l=0.5
X145 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=2 pd=14.7 as=2 ps=14.7 w=8 l=0.5
X146 cmfb_block_0/VREF cmfb_block_0/VREF VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.13 as=0.143 ps=1.06 w=0.5 l=0.5
X147 VOUT m1_6795_368# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.571 ps=4.24 w=2 l=0.5
C0 VCC folded_cascode_0/Vb2 3.37f
C1 VCC current_source_0/a_798_3689# 4.99f
C2 cmfb_block_0/a_2761_n1936# VCC 2.35f
C3 cmfb_block_0/IN cmfb_block_0/IP 1.42f
C4 input_stage_0/N2 input_stage_0/m1_n402_n3947# 1.63f
C5 current_source_0/li_226_2694# current_source_0/m1_1913_2070# 1.37f
C6 current_source_0/li_226_2694# current_source_0/li_805_1641# 1.31f
C7 VCC folded_cascode_0/Vb3 1.33f
C8 VCC cmfb_block_0/Vb1 6.27f
C9 input_stage_0/N3 input_stage_0/N4 3.91f
C10 cmfb_block_0/Vb1 folded_cascode_0/Vb2 1.22f
C11 cmfb_block_0/m1_3637_198# cmfb_block_0/CMFB 1.67f
C12 VSS cmfb_block_0/CMFB 5.99f
C13 input_stage_0/m1_n402_n3947# input_stage_0/N1 1.74f
C14 current_source_0/li_226_2694# current_source_0/li_1085_2889# 2.69f
C15 cmfb_block_0/IP VCC 1.5f
C16 VCC input_stage_0/N2 1.06f
C17 cmfb_block_0/VREF VCC 2.11f
C18 current_source_0/li_805_1641# folded_cascode_0/Vb2 1.06f
C19 VSS input_stage_0/m1_n402_n3947# 2.28f
C20 input_stage_0/m1_n402_90# input_stage_0/N4 1.63f
C21 current_source_0/m1_737_1534# current_source_0/li_805_1641# 1.06f
C22 VCC current_source_0/li_1085_2889# 2.04f
C23 VCC input_stage_0/N1 1.41f
C24 current_source_0/li_1085_2889# current_source_0/a_798_3689# 1.38f
C25 VCC VSS 2.54f
C26 input_stage_0/m1_n402_90# input_stage_0/N3 1.75f
C27 VCC input_stage_0/N3 1.09f
C28 input_stage_0/Vb5 VSS 3.89f
C29 current_source_0/li_1085_2889# folded_cascode_0/Vb3 1.01f
C30 current_source_0/li_1035_74# VSS 1.94f
C31 current_source_0/m1_1325_3826# VCC 1.51f
C32 VSS current_source_0/m1_737_1534# 2.37f
C33 cmfb_block_0/IN VCC 1.1f
C34 VCC current_source_0/li_226_2694# 1.15f
C35 cmfb_block_0/m1_3052_n816# cmfb_block_0/CMFB 1.95f
C36 current_source_0/li_226_2694# folded_cascode_0/Vb2 1.05f
C37 VCC diff_to_single_ended_1/a_n296_n44# 1.51f
C38 input_stage_0/N2 input_stage_0/N1 3.81f
C39 VCC input_stage_0/m1_n402_90# 3.03f
C40 VCC current_source_0/m1_737_3994# 2.41f
C41 VSS current_source_0/li_805_1641# 1.99f
C42 current_source_0/a_798_3689# current_source_0/m1_737_3994# 1.03f
C43 m1_6795_368# 0 1.05f
C44 input_stage_0/Vb5 0 3.91f
C45 cmfb_block_0/IN 0 1.56f
C46 input_stage_0/N1 0 1.52f
C47 cmfb_block_0/IP 0 1.52f
C48 input_stage_0/N2 0 1.74f
C49 input_stage_0/N3 0 1.16f
C50 diff_to_single_ended_1/a_n296_n44# 0 1.09f
C51 VOUT 0 1.18f
C52 cmfb_block_0/CMFB 0 3.31f
C53 cmfb_block_0/a_2761_n1936# 0 1.26f
C54 cmfb_block_0/VREF 0 1.79f
C55 current_source_0/li_226_2694# 0 5f
C56 cmfb_block_0/Vb1 0 1.61f
C57 VCC 0 82.1f
C58 current_source_0/a_798_3689# 0 3.2f
C59 current_source_0/m1_151_2991# 0 1.01f
C60 VSS 0 14.5f
C61 current_source_0/li_805_1641# 0 5.27f
C62 folded_cascode_0/Vb2 0 1.37f
C63 folded_cascode_0/Vb3 0 1.99f
C64 current_source_0/li_1085_2889# 0 2.34f
C65 current_source_0/li_1035_74# 0 1.8f
.ends
