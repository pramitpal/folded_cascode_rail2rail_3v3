** sch_path: /foss/designs/Comparator/old/schematic/folded_cascode/input_stage.sch
.subckt input_stage INN INP Vb1 Vb5 N1 N2 N3 N4 VCC VSS
*.PININFO INN:I INP:I Vb1:I Vb5:I N1:O N2:O N3:O N4:O VCC:I VSS:I
XM16 N2 INN net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM17 N1 INP net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM6 N3 INP net2 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM21 net2 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=4
XM18 net1 Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=4
XM4 N4 INN net2 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM2 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM3 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM5 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM7 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
XM8 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
XM9 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
XM10 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
.ends
.end
