magic
tech sky130A
magscale 1 2
timestamp 1696699629
<< mvnmos >>
rect -100 -81 100 19
<< mvndiff >>
rect -158 7 -100 19
rect -158 -69 -146 7
rect -112 -69 -100 7
rect -158 -81 -100 -69
rect 100 7 158 19
rect 100 -69 112 7
rect 146 -69 158 7
rect 100 -81 158 -69
<< mvndiffc >>
rect -146 -69 -112 7
rect 112 -69 146 7
<< poly >>
rect -100 91 100 107
rect -100 57 -84 91
rect 84 57 100 91
rect -100 19 100 57
rect -100 -107 100 -81
<< polycont >>
rect -84 57 84 91
<< locali >>
rect -100 57 -84 91
rect 84 57 100 91
rect -146 7 -112 23
rect -146 -85 -112 -69
rect 112 7 146 23
rect 112 -85 146 -69
<< viali >>
rect -84 57 84 91
rect -146 -69 -112 7
rect 112 -69 146 7
<< metal1 >>
rect -96 91 96 97
rect -96 57 -84 91
rect 84 57 96 91
rect -96 51 96 57
rect -152 7 -106 19
rect -152 -69 -146 7
rect -112 -69 -106 7
rect -152 -81 -106 -69
rect 106 7 152 19
rect 106 -69 112 7
rect 146 -69 152 7
rect 106 -81 152 -69
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
