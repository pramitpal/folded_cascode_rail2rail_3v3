magic
tech sky130A
magscale 1 2
timestamp 1697286120
<< nwell >>
rect 588 3022 6914 4593
rect 4105 2340 6914 3022
rect 4105 2117 6515 2340
rect 6106 1264 6911 1698
rect 6560 491 6908 1264
<< poly >>
rect 6684 2362 6784 2409
rect 6684 2328 6700 2362
rect 6768 2328 6784 2362
rect 6684 2312 6784 2328
rect 6684 2253 6784 2269
rect 6684 2219 6700 2253
rect 6768 2219 6784 2253
rect 6684 2172 6784 2219
rect 6684 415 6784 527
<< polycont >>
rect 6700 2328 6768 2362
rect 6700 2219 6768 2253
<< locali >>
rect 1785 4207 2263 4428
rect 329 4160 663 4194
rect 1222 4160 1585 4194
rect 1872 3832 1947 3866
rect 3410 3560 3752 3594
rect 3959 3131 4251 4351
rect 4853 4260 5058 4294
rect 5274 3177 6192 3211
rect 3828 2935 3976 2969
rect 2273 2856 2847 2890
rect 6340 2434 6658 4391
rect 6263 2421 6658 2434
rect -50 2187 -16 2275
rect -50 2153 23 2187
rect 1985 2065 2019 2373
rect 6263 2373 6482 2421
rect 2160 2065 2194 2373
rect 6261 2233 6482 2373
rect 6684 2328 6700 2362
rect 6768 2328 6784 2362
rect 6700 2310 6768 2328
rect 6700 2270 6713 2310
rect 6747 2270 6768 2310
rect 6700 2253 6768 2270
rect 2077 2031 2194 2065
rect 2077 261 2111 2031
rect 3926 1821 4234 2030
rect 3994 1820 4230 1821
rect 5276 1699 5310 1893
rect 6406 1582 6482 2233
rect 6684 2219 6700 2253
rect 6768 2219 6784 2253
rect 6406 1523 6647 1582
rect 6350 1447 6647 1523
rect 6431 1338 6647 1447
rect 5293 453 5327 492
rect 6356 327 6673 403
rect 1992 227 2111 261
rect 385 174 419 199
rect 5239 223 5344 271
rect 5239 175 5269 223
rect 5317 175 5344 223
rect 385 140 677 174
rect 5239 88 5344 175
rect 1797 28 1852 88
rect 1912 28 1914 88
rect 4216 82 5344 88
rect 4216 34 4222 82
rect 4270 34 5344 82
rect 4216 28 5344 34
<< viali >>
rect 295 4160 329 4194
rect 1585 4160 1619 4194
rect 1947 3832 1981 3866
rect 3752 3560 3786 3594
rect 4819 4260 4853 4294
rect 6192 3177 6226 3211
rect 3976 2932 4010 2972
rect 2239 2856 2273 2890
rect 1985 2373 2019 2407
rect 2160 2373 2194 2407
rect 6713 2270 6747 2310
rect 1985 2031 2019 2065
rect 6316 1844 6352 2006
rect 5276 1665 5310 1699
rect 5293 492 5327 526
rect 385 199 419 233
rect 1958 227 1992 261
rect 5269 175 5317 223
rect 1852 28 1912 88
rect 4222 34 4270 82
<< metal1 >>
rect 4118 4303 4170 4309
rect 4813 4303 4859 4306
rect 4046 4260 4118 4294
rect 289 4194 335 4206
rect -44 4160 295 4194
rect 329 4160 335 4194
rect 289 4148 335 4160
rect 1579 4194 1625 4206
rect 1579 4160 1585 4194
rect 1619 4160 2061 4194
rect 1579 4148 1625 4160
rect 1872 2292 1906 3921
rect 1938 3875 1990 3881
rect 1935 3826 1938 3872
rect 1990 3826 1993 3872
rect 1938 3817 1990 3823
rect 2027 3594 2061 4160
rect 3746 3594 3792 3606
rect 4046 3594 4080 4260
rect 4804 4251 4810 4303
rect 4862 4251 4868 4303
rect 4118 4245 4170 4251
rect 4813 4248 4859 4251
rect 2027 3560 2206 3594
rect 3746 3560 3752 3594
rect 3786 3560 4080 3594
rect 3746 3548 3792 3560
rect 2077 3417 2191 3451
rect 1979 2407 2025 2419
rect 2077 2407 2111 3417
rect 6186 3211 6232 3223
rect 6438 3211 6444 3220
rect 6186 3177 6192 3211
rect 6226 3177 6444 3211
rect 6186 3165 6232 3177
rect 6438 3168 6444 3177
rect 6496 3168 6502 3220
rect 3970 2978 4022 2984
rect 3964 2926 3970 2978
rect 3970 2920 4022 2926
rect 2233 2899 2279 2902
rect 2224 2847 2230 2899
rect 2282 2847 2288 2899
rect 2233 2844 2279 2847
rect 2154 2416 2200 2419
rect 1979 2373 1985 2407
rect 2019 2373 2111 2407
rect 1979 2361 2025 2373
rect 2145 2364 2151 2416
rect 2203 2364 2209 2416
rect 2154 2361 2200 2364
rect 6707 2316 6759 2322
rect 1872 2258 2607 2292
rect 6701 2264 6707 2316
rect 6707 2258 6759 2264
rect 6796 2304 6830 2479
rect 6865 2304 6871 2313
rect 6796 2270 6871 2304
rect -50 2153 50 2187
rect -50 2076 -16 2153
rect 1979 2065 2025 2077
rect 1979 2031 1985 2065
rect 2019 2031 2111 2065
rect 1979 2019 2025 2031
rect 2077 270 2111 2031
rect 4064 1795 4098 2201
rect 6310 2006 6667 2030
rect 4752 1795 4758 1804
rect 4064 1761 4758 1795
rect 4752 1752 4758 1761
rect 4810 1795 4816 1804
rect 5276 1795 5310 1865
rect 6310 1844 6316 2006
rect 6352 1958 6667 2006
rect 6352 1844 6669 1958
rect 6310 1820 6669 1844
rect 4810 1761 5310 1795
rect 6796 1784 6830 2270
rect 6865 2261 6871 2270
rect 6923 2261 6929 2313
rect 4810 1752 4816 1761
rect 5267 1708 5319 1714
rect 5264 1659 5267 1705
rect 5319 1659 5322 1705
rect 5267 1650 5319 1656
rect 6781 1653 6787 1705
rect 6839 1653 6845 1705
rect 6796 1568 6830 1653
rect 4130 1377 4136 1429
rect 4188 1377 4194 1429
rect 4145 1276 4179 1377
rect 4145 1242 4230 1276
rect 6804 612 6901 646
rect 6496 553 6548 559
rect 5284 535 5336 541
rect 5281 486 5284 532
rect 5336 486 5339 532
rect 6548 510 6726 544
rect 6496 495 6548 501
rect 5284 477 5336 483
rect 6867 402 6901 612
rect 6795 368 6901 402
rect 1946 261 2004 267
rect 376 242 428 248
rect 373 193 376 239
rect 428 193 431 239
rect 1946 227 1958 261
rect 1992 227 2004 261
rect 1946 221 2004 227
rect 2062 218 2068 270
rect 2120 218 2126 270
rect 5263 229 5323 235
rect 376 184 428 190
rect 5257 169 5263 229
rect 5323 169 5329 229
rect 5263 163 5323 169
rect 1846 94 1918 100
rect 1846 88 1858 94
rect 1846 28 1852 88
rect 1846 22 1858 28
rect 1918 22 1924 94
rect 4216 88 4276 94
rect 4210 28 4216 88
rect 4276 28 4282 88
rect 4216 22 4276 28
rect 1846 16 1918 22
<< via1 >>
rect 1938 3866 1990 3875
rect 1938 3832 1947 3866
rect 1947 3832 1981 3866
rect 1981 3832 1990 3866
rect 1938 3823 1990 3832
rect 4118 4251 4170 4303
rect 4810 4294 4862 4303
rect 4810 4260 4819 4294
rect 4819 4260 4853 4294
rect 4853 4260 4862 4294
rect 4810 4251 4862 4260
rect 6444 3168 6496 3220
rect 3970 2972 4022 2978
rect 3970 2932 3976 2972
rect 3976 2932 4010 2972
rect 4010 2932 4022 2972
rect 3970 2926 4022 2932
rect 2230 2890 2282 2899
rect 2230 2856 2239 2890
rect 2239 2856 2273 2890
rect 2273 2856 2282 2890
rect 2230 2847 2282 2856
rect 2151 2407 2203 2416
rect 2151 2373 2160 2407
rect 2160 2373 2194 2407
rect 2194 2373 2203 2407
rect 2151 2364 2203 2373
rect 6707 2310 6759 2316
rect 6707 2270 6713 2310
rect 6713 2270 6747 2310
rect 6747 2270 6759 2310
rect 6707 2264 6759 2270
rect 4758 1752 4810 1804
rect 6871 2261 6923 2313
rect 5267 1699 5319 1708
rect 5267 1665 5276 1699
rect 5276 1665 5310 1699
rect 5310 1665 5319 1699
rect 5267 1656 5319 1665
rect 6787 1653 6839 1705
rect 4136 1377 4188 1429
rect 5284 526 5336 535
rect 5284 492 5293 526
rect 5293 492 5327 526
rect 5327 492 5336 526
rect 5284 483 5336 492
rect 6496 501 6548 553
rect 376 233 428 242
rect 376 199 385 233
rect 385 199 419 233
rect 419 199 428 233
rect 376 190 428 199
rect 2068 218 2120 270
rect 5263 223 5323 229
rect 5263 175 5269 223
rect 5269 175 5317 223
rect 5317 175 5323 223
rect 5263 169 5323 175
rect 1858 88 1918 94
rect 1858 28 1912 88
rect 1912 28 1918 88
rect 1858 22 1918 28
rect 4216 82 4276 88
rect 4216 34 4222 82
rect 4222 34 4270 82
rect 4270 34 4276 82
rect 4216 28 4276 34
<< metal2 >>
rect 4810 4303 4862 4309
rect 4112 4251 4118 4303
rect 4170 4294 4176 4303
rect 4170 4260 4810 4294
rect 4170 4251 4176 4260
rect 4810 4245 4862 4251
rect 1947 3875 1981 3882
rect 1932 3823 1938 3875
rect 1990 3823 1996 3875
rect 1554 3539 1610 3548
rect -44 3494 1554 3528
rect 1554 3474 1610 3483
rect 1557 2890 1566 2901
rect -117 2856 1566 2890
rect 1557 2845 1566 2856
rect 1622 2845 1631 2901
rect 1947 2292 1981 3823
rect 2035 3481 2044 3541
rect 2104 3528 2113 3541
rect 2104 3494 2191 3528
rect 2104 3481 2113 3494
rect 2077 3417 2449 3451
rect 2077 2407 2111 3417
rect 4132 3341 4192 3350
rect 4132 3272 4192 3281
rect 6444 3220 6496 3226
rect 6496 3177 6976 3211
rect 6444 3162 6496 3168
rect 3701 2922 3710 2982
rect 3770 2922 3779 2982
rect 3964 2926 3970 2978
rect 4022 2969 4028 2978
rect 4145 2969 4179 3090
rect 4022 2935 4179 2969
rect 4022 2926 4028 2935
rect 2230 2903 2282 2905
rect 2217 2843 2226 2903
rect 2286 2843 2295 2903
rect 2230 2841 2282 2843
rect 2151 2416 2203 2422
rect 2077 2373 2151 2407
rect 2151 2358 2203 2364
rect 1947 2258 2784 2292
rect 4145 1435 4179 2935
rect 6701 2264 6707 2316
rect 6759 2264 6765 2316
rect 6871 2313 6923 2319
rect 4758 1808 4810 1810
rect 4745 1748 4754 1808
rect 4814 1748 4823 1808
rect 4758 1746 4810 1748
rect 5261 1656 5267 1708
rect 5319 1656 5325 1708
rect 6716 1696 6750 2264
rect 6923 2270 6987 2304
rect 6871 2255 6923 2261
rect 6787 1705 6839 1711
rect 6716 1662 6787 1696
rect 4136 1429 4188 1435
rect 4136 1371 4188 1377
rect 4172 1171 4181 1231
rect 4241 1218 4250 1231
rect 4241 1184 4281 1218
rect 4241 1171 4250 1184
rect 5276 700 5310 1656
rect 6787 1647 6839 1653
rect 6273 1188 6539 1222
rect 5263 691 5323 700
rect 5263 622 5323 631
rect 6505 553 6539 1188
rect 5278 526 5284 535
rect -24 492 5284 526
rect 385 242 419 492
rect 5278 483 5284 492
rect 5336 483 5342 535
rect 6490 501 6496 553
rect 6548 501 6554 553
rect 2068 270 2120 276
rect 370 190 376 242
rect 428 190 434 242
rect 1890 227 2068 261
rect 5263 229 5323 235
rect 2068 212 2120 218
rect 5256 171 5263 227
rect 5323 171 5330 227
rect 5263 163 5323 169
rect 1858 94 1918 100
rect 1849 22 1858 94
rect 1918 22 1927 94
rect 4218 88 4274 95
rect 4210 28 4216 88
rect 4276 28 4282 88
rect 1858 16 1918 22
rect 4218 21 4274 28
<< via2 >>
rect 1554 3483 1610 3539
rect 1566 2845 1622 2901
rect 2044 3481 2104 3541
rect 4132 3281 4192 3341
rect 3710 2922 3770 2982
rect 2226 2899 2286 2903
rect 2226 2847 2230 2899
rect 2230 2847 2282 2899
rect 2282 2847 2286 2899
rect 2226 2843 2286 2847
rect 4754 1804 4814 1808
rect 4754 1752 4758 1804
rect 4758 1752 4810 1804
rect 4810 1752 4814 1804
rect 4754 1748 4814 1752
rect 4181 1171 4241 1231
rect 5263 631 5323 691
rect 5265 171 5321 227
rect 1858 22 1918 94
rect 4218 30 4274 86
<< metal3 >>
rect 1549 3541 1615 3544
rect 2039 3541 2109 3546
rect 1549 3539 2044 3541
rect 1549 3483 1554 3539
rect 1610 3483 2044 3539
rect 1549 3481 2044 3483
rect 2104 3481 2109 3541
rect 1549 3478 1615 3481
rect 2039 3476 2109 3481
rect 4127 3341 4197 3346
rect 4127 3281 4132 3341
rect 4192 3281 4197 3341
rect 4127 3276 4197 3281
rect 3705 2982 3775 2987
rect 4132 2982 4192 3276
rect 3705 2922 3710 2982
rect 3770 2922 4192 2982
rect 3705 2917 3775 2922
rect 1561 2903 1627 2906
rect 2221 2903 2291 2908
rect 1561 2901 2226 2903
rect 1561 2845 1566 2901
rect 1622 2845 2226 2901
rect 1561 2843 2226 2845
rect 2286 2843 2291 2903
rect 1561 2840 1627 2843
rect 2221 2838 2291 2843
rect 4048 1231 4108 2922
rect 4294 1746 4300 1810
rect 4364 1808 4370 1810
rect 4749 1808 4819 1813
rect 4364 1748 4754 1808
rect 4814 1748 4819 1808
rect 4364 1746 4370 1748
rect 4749 1743 4819 1748
rect 4176 1231 4246 1236
rect 4048 1171 4181 1231
rect 4241 1171 4246 1231
rect 4176 1166 4246 1171
rect 5258 691 5328 696
rect 5258 631 5263 691
rect 5323 631 5328 691
rect 5258 626 5328 631
rect 5263 232 5323 626
rect 5260 227 5326 232
rect 5260 171 5265 227
rect 5321 171 5326 227
rect 5260 166 5326 171
rect 1853 94 1923 99
rect 1853 22 1858 94
rect 1918 88 1923 94
rect 4213 88 4279 91
rect 1918 86 4279 88
rect 1918 30 4218 86
rect 4274 30 4279 86
rect 1918 28 4279 30
rect 1918 22 1923 28
rect 4213 25 4279 28
rect 1853 17 1923 22
<< via3 >>
rect 4300 1746 4364 1810
<< metal4 >>
rect 4299 1810 4365 1811
rect 4299 1808 4300 1810
rect 3164 1748 4300 1808
rect 3164 998 3224 1748
rect 4299 1746 4300 1748
rect 4364 1746 4365 1810
rect 4299 1745 4365 1746
use cmfb_block  cmfb_block_0 /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/layout/cmfb
timestamp 1697281155
transform 1 0 1927 0 1 3940
box 2178 -2124 4555 634
use diff_to_single_ended  diff_to_single_ended_1 /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/layout/diff_to_single_ended
timestamp 1697284980
transform 1 0 4992 0 1 1355
box -906 -1112 1548 343
use folded_cascode  folded_cascode_0 /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/layout/folded_cascode
timestamp 1697281155
transform 1 0 2899 0 1 3365
box -742 -2133 1199 1176
use input_stage  input_stage_0 /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/layout/input_stage
timestamp 1697284980
transform 1 0 890 0 1 4022
box -901 -4108 1102 571
use sky130_fd_pr__cap_mim_m3_1_N2QRHY  sky130_fd_pr__cap_mim_m3_1_N2QRHY_0
timestamp 1697281155
transform 1 0 3070 0 1 588
box -896 -640 896 640
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_0 /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/layout/diff_to_single_ended
timestamp 1697284980
transform 1 0 6734 0 1 1972
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_VNB5GC  sky130_fd_pr__nfet_g5v0d10v5_VNB5GC_0 /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/layout/diff_to_single_ended
timestamp 1697284980
transform 1 0 6734 0 1 365
box -108 -76 108 76
use sky130_fd_pr__pfet_g5v0d10v5_2V6JZ7  sky130_fd_pr__pfet_g5v0d10v5_2V6JZ7_0
timestamp 1697286120
transform 1 0 6734 0 1 3409
box -174 -1066 174 1066
use sky130_fd_pr__pfet_g5v0d10v5_GX3LZ5  sky130_fd_pr__pfet_g5v0d10v5_GX3LZ5_0
timestamp 1697286120
transform 1 0 6734 0 1 1055
box -174 -564 174 602
<< labels >>
flabel metal1 s -34 4175 -34 4175 0 FreeSans 800 0 0 0 Vb1
flabel metal2 s -30 3515 -30 3515 0 FreeSans 800 0 0 0 Vb2
flabel metal2 s -105 2872 -105 2872 0 FreeSans 800 0 0 0 Vb3
flabel metal2 s -11 509 -11 509 0 FreeSans 800 0 0 0 Vb5
flabel locali s 2021 4344 2021 4344 0 FreeSans 800 0 0 0 VCC
flabel locali s 5296 84 5296 84 0 FreeSans 800 0 0 0 VSS
flabel metal1 s -36 2090 -36 2090 0 FreeSans 800 0 0 0 INP
flabel locali s -35 2262 -35 2262 0 FreeSans 800 0 0 0 INN
flabel metal2 s 6519 1206 6519 1206 0 FreeSans 800 0 0 0 V
flabel metal2 s 6971 2288 6971 2288 0 FreeSans 800 0 0 0 VOUT
flabel metal2 s 6961 3196 6961 3196 0 FreeSans 800 0 0 0 VREF
<< end >>
