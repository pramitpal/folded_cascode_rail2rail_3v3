magic
tech sky130A
magscale 1 2
timestamp 1697289488
<< error_p >>
rect -144 80 144 114
rect -174 -152 174 80
<< nwell >>
rect -144 -148 144 114
<< mvpmos >>
rect -50 -86 50 14
<< mvpdiff >>
rect -108 2 -50 14
rect -108 -74 -96 2
rect -62 -74 -50 2
rect -108 -86 -50 -74
rect 50 2 108 14
rect 50 -74 62 2
rect 96 -74 108 2
rect 50 -86 108 -74
<< mvpdiffc >>
rect -96 -74 -62 2
rect 62 -74 96 2
<< poly >>
rect -50 95 50 111
rect -50 61 -34 95
rect 34 61 50 95
rect -50 14 50 61
rect -50 -112 50 -86
<< polycont >>
rect -34 61 34 95
<< locali >>
rect -50 61 -34 95
rect 34 61 50 95
rect -96 2 -62 18
rect -96 -90 -62 -74
rect 62 2 96 18
rect 62 -90 96 -74
<< viali >>
rect -34 61 34 95
rect -96 -74 -62 2
rect 62 -74 96 2
<< metal1 >>
rect -46 95 46 101
rect -46 61 -34 95
rect 34 61 46 95
rect -46 55 46 61
rect -102 2 -56 14
rect -102 -74 -96 2
rect -62 -74 -56 2
rect -102 -86 -56 -74
rect 56 2 102 14
rect 56 -74 62 2
rect 96 -74 102 2
rect 56 -86 102 -74
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
