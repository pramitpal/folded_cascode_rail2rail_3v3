magic
tech sky130A
magscale 1 2
timestamp 1698929273
<< error_p >>
rect -258 -331 -200 269
rect 200 -331 258 269
<< mvnmos >>
rect -200 -331 200 269
<< mvndiff >>
rect -258 257 -200 269
rect -258 -319 -246 257
rect -212 -319 -200 257
rect -258 -331 -200 -319
rect 200 257 258 269
rect 200 -319 212 257
rect 246 -319 258 257
rect 200 -331 258 -319
<< mvndiffc >>
rect -246 -319 -212 257
rect 212 -319 246 257
<< poly >>
rect -200 341 200 357
rect -200 307 -184 341
rect 184 307 200 341
rect -200 269 200 307
rect -200 -357 200 -331
<< polycont >>
rect -184 307 184 341
<< locali >>
rect -200 307 -184 341
rect 184 307 200 341
rect -246 257 -212 273
rect -246 -335 -212 -319
rect 212 257 246 273
rect 212 -335 246 -319
<< viali >>
rect -184 307 184 341
rect -246 -319 -212 257
rect 212 -319 246 257
<< metal1 >>
rect -196 341 196 347
rect -196 307 -184 341
rect 184 307 196 341
rect -196 301 196 307
rect -252 257 -206 269
rect -252 -319 -246 257
rect -212 -319 -206 257
rect -252 -331 -206 -319
rect 206 257 252 269
rect 206 -319 212 257
rect 246 -319 252 257
rect 206 -331 252 -319
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
