magic
tech sky130A
magscale 1 2
timestamp 1698929273
<< error_p >>
rect -258 -431 -200 369
rect 200 -431 258 369
<< mvnmos >>
rect -200 -431 200 369
<< mvndiff >>
rect -258 357 -200 369
rect -258 -419 -246 357
rect -212 -419 -200 357
rect -258 -431 -200 -419
rect 200 357 258 369
rect 200 -419 212 357
rect 246 -419 258 357
rect 200 -431 258 -419
<< mvndiffc >>
rect -246 -419 -212 357
rect 212 -419 246 357
<< poly >>
rect -200 441 200 457
rect -200 407 -184 441
rect 184 407 200 441
rect -200 369 200 407
rect -200 -457 200 -431
<< polycont >>
rect -184 407 184 441
<< locali >>
rect -200 407 -184 441
rect 184 407 200 441
rect -246 357 -212 373
rect -246 -435 -212 -419
rect 212 357 246 373
rect 212 -435 246 -419
<< viali >>
rect -184 407 184 441
rect -246 -419 -212 357
rect 212 -419 246 357
<< metal1 >>
rect -196 441 196 447
rect -196 407 -184 441
rect 184 407 196 441
rect -196 401 196 407
rect -252 357 -206 369
rect -252 -419 -246 357
rect -212 -419 -206 357
rect -252 -431 -206 -419
rect 206 357 252 369
rect 206 -419 212 357
rect 246 -419 252 357
rect 206 -431 252 -419
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
