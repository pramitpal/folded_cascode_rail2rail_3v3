magic
tech sky130A
magscale 1 2
timestamp 1696699961
<< mvnmos >>
rect -250 -81 250 19
<< mvndiff >>
rect -308 7 -250 19
rect -308 -69 -296 7
rect -262 -69 -250 7
rect -308 -81 -250 -69
rect 250 7 308 19
rect 250 -69 262 7
rect 296 -69 308 7
rect 250 -81 308 -69
<< mvndiffc >>
rect -296 -69 -262 7
rect 262 -69 296 7
<< poly >>
rect -250 91 250 107
rect -250 57 -234 91
rect 234 57 250 91
rect -250 19 250 57
rect -250 -107 250 -81
<< polycont >>
rect -234 57 234 91
<< locali >>
rect -250 57 -234 91
rect 234 57 250 91
rect -296 7 -262 23
rect -296 -85 -262 -69
rect 262 7 296 23
rect 262 -85 296 -69
<< viali >>
rect -234 57 234 91
rect -296 -69 -262 7
rect 262 -69 296 7
<< metal1 >>
rect -246 91 246 97
rect -246 57 -234 91
rect 234 57 246 91
rect -246 51 246 57
rect -302 7 -256 19
rect -302 -69 -296 7
rect -262 -69 -256 7
rect -302 -81 -256 -69
rect 256 7 302 19
rect 256 -69 262 7
rect 296 -69 302 7
rect 256 -81 302 -69
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 2.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
