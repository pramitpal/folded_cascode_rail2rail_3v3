magic
tech sky130A
magscale 1 2
timestamp 1698920341
<< mvnmos >>
rect -50 -1331 50 1269
<< mvndiff >>
rect -108 1257 -50 1269
rect -108 -1319 -96 1257
rect -62 -1319 -50 1257
rect -108 -1331 -50 -1319
rect 50 1257 108 1269
rect 50 -1319 62 1257
rect 96 -1319 108 1257
rect 50 -1331 108 -1319
<< mvndiffc >>
rect -96 -1319 -62 1257
rect 62 -1319 96 1257
<< poly >>
rect -50 1341 50 1357
rect -50 1307 -34 1341
rect 34 1307 50 1341
rect -50 1269 50 1307
rect -50 -1357 50 -1331
<< polycont >>
rect -34 1307 34 1341
<< locali >>
rect -50 1307 -34 1341
rect 34 1307 50 1341
rect -96 1257 -62 1273
rect -96 -1335 -62 -1319
rect 62 1257 96 1273
rect 62 -1335 96 -1319
<< viali >>
rect -34 1307 34 1341
rect -96 -1319 -62 1257
rect 62 -1319 96 1257
<< metal1 >>
rect -46 1341 46 1347
rect -46 1307 -34 1341
rect 34 1307 46 1341
rect -46 1301 46 1307
rect -102 1257 -56 1269
rect -102 -1319 -96 1257
rect -62 -1319 -56 1257
rect -102 -1331 -56 -1319
rect 56 1257 102 1269
rect 56 -1319 62 1257
rect 96 -1319 102 1257
rect 56 -1331 102 -1319
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 13 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
