* NGSPICE file created from total.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_VNB5GC a_n108_n50# a_50_n50# a_n50_n76# VSUBS
X0 a_50_n50# a_n50_n76# a_n108_n50# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__res_generic_nd__hv_USEA7F a_n114_n346# a_30_n346# VSUBS
X0 a_30_n346# a_n114_n346# VSUBS sky130_fd_pr__res_generic_nd__hv w=0.415 l=5.8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_MBRSZA a_n258_n264# a_n200_n361# a_200_n264#
+ w_n294_n364#
X0 a_200_n264# a_n200_n361# a_n258_n264# w_n294_n364# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_EHRSHC a_n258_n400# w_n294_n462# a_200_n400#
+ a_n200_n426#
X0 a_200_n400# a_n200_n426# a_n258_n400# w_n294_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_K5LT42 a_n258_n331# a_200_n331# a_n200_n357#
+ VSUBS
X0 a_200_n331# a_n200_n357# a_n258_n331# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NYRQZ6 a_n108_n231# a_50_n231# a_n50_n257# VSUBS
X0 a_50_n231# a_n50_n257# a_n108_n231# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CMVU23 a_200_n831# a_n200_n857# a_n258_n831#
+ VSUBS
X0 a_200_n831# a_n200_n857# a_n258_n831# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CM22X2 a_200_n431# a_n200_n457# a_n258_n431#
+ VSUBS
X0 a_200_n431# a_n200_n457# a_n258_n431# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TNTUPH a_50_n431# a_n50_n457# a_n108_n431# VSUBS
X0 a_50_n431# a_n50_n457# a_n108_n431# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_JSTQTR a_50_n1351# a_n50_n1377# a_n108_n1351#
+ VSUBS
X0 a_50_n1351# a_n50_n1377# a_n108_n1351# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=3.83 pd=27 as=3.83 ps=27 w=13.2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5 a_n108_n764# a_n50_n861# a_50_n764# w_n144_n864#
X0 a_50_n764# a_n50_n861# a_n108_n764# w_n144_n864# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_KRRUZH a_n50_n597# a_n108_n571# a_50_n571# VSUBS
X0 a_50_n571# a_n50_n597# a_n108_n571# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.57 pd=11.4 as=1.57 ps=11.4 w=5.4 l=0.5
.ends

.subckt current_source Vb5 VSS Vb3 Vb2 Vb1 VCC
Xsky130_fd_pr__res_generic_nd__hv_USEA7F_2 li_1035_74# VSS VSS sky130_fd_pr__res_generic_nd__hv_USEA7F
Xsky130_fd_pr__res_generic_nd__hv_USEA7F_3 VSS li_1035_74# VSS sky130_fd_pr__res_generic_nd__hv_USEA7F
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_6 m1_737_3994# li_1085_2889# Vb3 VCC sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_7 m1_1325_3826# li_1085_2889# li_226_2694# VCC
+ sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_2 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_8 Vb3 li_1085_2889# m1_737_3994# VCC sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_9 li_226_2694# li_1085_2889# m1_1325_3826# VCC
+ sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_3 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__nfet_g5v0d10v5_K5LT42_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_K5LT42
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_6 m1_737_3994# VCC VCC a_798_3689# sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__nfet_g5v0d10v5_NYRQZ6_0 Vb3 Vb5 Vb3 VSS sky130_fd_pr__nfet_g5v0d10v5_NYRQZ6
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_7 m1_1325_3826# VCC VCC a_798_3689# sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_8 a_798_3689# VCC VCC a_798_3689# sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_9 VCC VCC a_798_3689# a_798_3689# sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__nfet_g5v0d10v5_CMVU23_0 m1_1913_2070# li_805_1641# li_1035_74# VSS
+ sky130_fd_pr__nfet_g5v0d10v5_CMVU23
Xsky130_fd_pr__nfet_g5v0d10v5_CMVU23_2 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CMVU23
Xsky130_fd_pr__nfet_g5v0d10v5_CMVU23_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CMVU23
Xsky130_fd_pr__nfet_g5v0d10v5_CMVU23_3 li_1035_74# li_805_1641# m1_1913_2070# VSS
+ sky130_fd_pr__nfet_g5v0d10v5_CMVU23
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_10 a_798_3689# li_1085_2889# li_1085_2889# VCC
+ sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_11 li_1085_2889# li_1085_2889# a_798_3689# VCC
+ sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_0 Vb2 li_226_2694# m1_737_1534# VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_1 li_226_2694# li_226_2694# li_805_1641# VSS
+ sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_2 li_1085_2889# li_226_2694# m1_1913_2070# VSS
+ sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_TNTUPH_1 Vb5 Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5_TNTUPH
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_3 m1_1913_2070# li_226_2694# li_1085_2889# VSS
+ sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_10 VCC VCC m1_1325_3826# a_798_3689# sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_4 li_805_1641# li_226_2694# li_226_2694# VSS
+ sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_5 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__pfet_g5v0d10v5_EHRSHC_11 VCC VCC m1_737_3994# a_798_3689# sky130_fd_pr__pfet_g5v0d10v5_EHRSHC
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_6 li_805_1641# li_805_1641# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_7 VSS li_805_1641# li_805_1641# VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_10 VSS li_805_1641# m1_737_1534# VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_8 m1_737_1534# li_805_1641# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_11 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_JSTQTR_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_JSTQTR
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_12 m1_737_1534# li_226_2694# Vb2 VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_9 VSS m1_151_2991# a_798_3689# VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_JSTQTR_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_JSTQTR
Xsky130_fd_pr__nfet_g5v0d10v5_CM22X2_13 VSS li_226_2694# m1_151_2991# VSS sky130_fd_pr__nfet_g5v0d10v5_CM22X2
Xsky130_fd_pr__nfet_g5v0d10v5_JSTQTR_2 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_JSTQTR
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_0 Vb1 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5
Xsky130_fd_pr__nfet_g5v0d10v5_KRRUZH_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_KRRUZH
Xsky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_2 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_2 Vb2 Vb2 Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5
Xsky130_fd_pr__res_generic_nd__hv_USEA7F_0 li_1035_74# VSS VSS sky130_fd_pr__res_generic_nd__hv_USEA7F
Xsky130_fd_pr__pfet_g5v0d10v5_MBRSZA_3 m1_151_2991# li_226_2694# VCC VCC sky130_fd_pr__pfet_g5v0d10v5_MBRSZA
Xsky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_3 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5
Xsky130_fd_pr__res_generic_nd__hv_USEA7F_1 VSS li_1035_74# VSS sky130_fd_pr__res_generic_nd__hv_USEA7F
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_JEERZ7 w_n144_n462# a_50_n400# a_n50_n426# a_n108_n400#
X0 a_50_n400# a_n50_n426# a_n108_n400# w_n144_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6LM9S7 a_n108_n50# w_n144_n112# a_50_n50# a_n50_n76#
X0 a_50_n50# a_n50_n76# a_n108_n50# w_n144_n112# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7JP9SF a_n208_n86# a_150_n86# a_n150_n112# w_n244_n148#
X0 a_150_n86# a_n150_n112# a_n208_n86# w_n244_n148# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_6DL6AA a_100_n50# a_n100_n76# a_n158_n50# VSUBS
X0 a_100_n50# a_n100_n76# a_n158_n50# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GUWUK4 a_n108_n19# a_n50_n107# a_50_n19# VSUBS
X0 a_50_n19# a_n50_n107# a_n108_n19# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3JERZF w_n244_n498# a_150_n436# a_n208_n436#
+ a_n150_n462#
X0 a_150_n436# a_n150_n462# a_n208_n436# w_n244_n498# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1.5
.ends

.subckt cmfb_block Vb1 CMFB VREF IP VCC VSS IN
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_10 VCC m1_3052_n816# VREF CMFB sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_11 VCC CMFB VREF m1_3052_n816# sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_12 VCC a_2761_n1936# IN m1_3637_198# sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__pfet_g5v0d10v5_6LM9S7_4 m1_3637_198# VCC VCC Vb1 sky130_fd_pr__pfet_g5v0d10v5_6LM9S7
Xsky130_fd_pr__pfet_g5v0d10v5_6LM9S7_5 VCC VCC m1_3052_n816# Vb1 sky130_fd_pr__pfet_g5v0d10v5_6LM9S7
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_13 VCC m1_3637_198# IN a_2761_n1936# sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__pfet_g5v0d10v5_6LM9S7_6 m1_3052_n816# VCC VCC Vb1 sky130_fd_pr__pfet_g5v0d10v5_6LM9S7
Xsky130_fd_pr__pfet_g5v0d10v5_7JP9SF_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_7JP9SF
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_14 VCC m1_3637_198# VREF CMFB sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__pfet_g5v0d10v5_7JP9SF_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_7JP9SF
Xsky130_fd_pr__pfet_g5v0d10v5_6LM9S7_7 VCC VCC m1_3637_198# Vb1 sky130_fd_pr__pfet_g5v0d10v5_6LM9S7
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_15 VCC CMFB VREF m1_3637_198# sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_8 VCC a_2761_n1936# IP m1_3052_n816# sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_9 VCC m1_3052_n816# IP a_2761_n1936# sky130_fd_pr__pfet_g5v0d10v5_JEERZ7
Xsky130_fd_pr__nfet_g5v0d10v5_6DL6AA_0 VSS CMFB CMFB VSS sky130_fd_pr__nfet_g5v0d10v5_6DL6AA
Xsky130_fd_pr__nfet_g5v0d10v5_GUWUK4_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_GUWUK4
Xsky130_fd_pr__nfet_g5v0d10v5_GUWUK4_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_GUWUK4
Xsky130_fd_pr__nfet_g5v0d10v5_6DL6AA_1 VSS a_2761_n1936# a_2761_n1936# VSS sky130_fd_pr__nfet_g5v0d10v5_6DL6AA
Xsky130_fd_pr__nfet_g5v0d10v5_6DL6AA_2 CMFB CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5_6DL6AA
Xsky130_fd_pr__nfet_g5v0d10v5_6DL6AA_3 a_2761_n1936# a_2761_n1936# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_6DL6AA
Xsky130_fd_pr__pfet_g5v0d10v5_3JERZF_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_3JERZF
Xsky130_fd_pr__pfet_g5v0d10v5_3JERZF_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_3JERZF
Xsky130_fd_pr__pfet_g5v0d10v5_3JERZF_2 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_3JERZF
Xsky130_fd_pr__pfet_g5v0d10v5_3JERZF_3 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_3JERZF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_N2QRHY m3_n896_n640# c1_n856_n600#
X0 c1_n856_n600# m3_n896_n640# sky130_fd_pr__cap_mim_m3_1 l=6 w=7.1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_2V6JZ7 a_n108_n1000# a_50_n1000# w_n144_n1062#
+ a_n50_n1026#
X0 a_50_n1000# a_n50_n1026# a_n108_n1000# w_n144_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_GX3LZ5 a_n108_n464# a_n50_n561# a_50_n464# w_n144_n564#
X0 a_50_n464# a_n50_n561# a_n108_n464# w_n144_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NY97Z6 a_50_n200# a_n50_n226# a_n108_n200# VSUBS
X0 a_50_n200# a_n50_n226# a_n108_n200# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CDSXD6 a_n258_n81# a_200_n81# a_n200_n107# VSUBS
X0 a_200_n81# a_n200_n107# a_n258_n81# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DFFFYB a_n200_n257# a_200_n169# a_n258_n169#
+ VSUBS
X0 a_200_n169# a_n200_n257# a_n258_n169# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HGG9EV a_100_n50# a_n100_n76# w_n194_n112# a_n158_n50#
X0 a_100_n50# a_n100_n76# a_n158_n50# w_n194_n112# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HCV9S7 a_n108_n86# w_n144_n148# a_50_n86# a_n50_n112#
X0 a_50_n86# a_n50_n112# a_n108_n86# w_n144_n148# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt diff_to_single_ended out vb5 v out2 VCC VSS
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_4 a_n296_n44# out li_n130_n833# VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_0 li_n130_n833# VSS vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_1 VSS li_n130_n833# vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC
Xsky130_fd_pr__nfet_g5v0d10v5_CDSXD6_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CDSXD6
Xsky130_fd_pr__nfet_g5v0d10v5_CDSXD6_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_CDSXD6
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_2 VSS li_n130_n833# vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_3 li_n130_n833# VSS vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC
Xsky130_fd_pr__nfet_g5v0d10v5_DFFFYB_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_DFFFYB
Xsky130_fd_pr__nfet_g5v0d10v5_DFFFYB_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_DFFFYB
Xsky130_fd_pr__pfet_g5v0d10v5_HGG9EV_0 VCC a_n296_n44# VCC a_n296_n44# sky130_fd_pr__pfet_g5v0d10v5_HGG9EV
Xsky130_fd_pr__pfet_g5v0d10v5_HGG9EV_2 v a_n296_n44# VCC VCC sky130_fd_pr__pfet_g5v0d10v5_HGG9EV
Xsky130_fd_pr__pfet_g5v0d10v5_HGG9EV_1 VCC a_n296_n44# VCC v sky130_fd_pr__pfet_g5v0d10v5_HGG9EV
Xsky130_fd_pr__pfet_g5v0d10v5_HGG9EV_3 a_n296_n44# a_n296_n44# VCC VCC sky130_fd_pr__pfet_g5v0d10v5_HGG9EV
Xsky130_fd_pr__pfet_g5v0d10v5_HCV9S7_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_HCV9S7
Xsky130_fd_pr__pfet_g5v0d10v5_HCV9S7_2 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_HCV9S7
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_0 li_n130_n833# out2 v VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_2 v out2 li_n130_n833# VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_3 li_n130_n833# out a_n296_n44# VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TNTUPH#0 a_50_n431# a_n50_n457# a_n108_n431#
+ VSUBS
X0 a_50_n431# a_n50_n457# a_n108_n431# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0 w_n144_n462# a_50_n400# a_n50_n426#
+ a_n108_n400#
X0 a_50_n400# a_n50_n426# a_n108_n400# w_n144_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0 a_50_n200# a_n50_n226# a_n108_n200#
+ VSUBS
X0 a_50_n200# a_n50_n226# a_n108_n200# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TNBBPH a_50_n400# a_n50_n426# a_n108_n400# VSUBS
X0 a_50_n400# a_n50_n426# a_n108_n400# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TNWANH a_n50_n457# a_50_n369# a_n108_n369# VSUBS
X0 a_50_n369# a_n50_n457# a_n108_n369# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7 w_n144_n162# a_50_n100# a_n50_n126# a_n108_n100#
X0 a_50_n100# a_n50_n126# a_n108_n100# w_n144_n162# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NYY6SB a_50_n169# a_n108_n169# a_n50_n257# VSUBS
X0 a_50_n169# a_n50_n257# a_n108_n169# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7 a_50_n136# a_n108_n136# a_n50_n162# w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_DEERZ7 a_50_n436# a_n108_n436# a_n50_n462# w_n144_n498#
X0 a_50_n436# a_n50_n462# a_n108_n436# w_n144_n498# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt folded_cascode Vb3 Vb2 Vb1 CMFB out N4 N3 N2 out2 N1 VCC VSS
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_2 VCC N2 Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_1 VCC VCC Vb1 N2 sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_4 N3 Vb3 out2 VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0
Xsky130_fd_pr__nfet_g5v0d10v5_TNBBPH_0 N3 CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5_TNBBPH
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_3 VCC VCC Vb1 N1 sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0
Xsky130_fd_pr__nfet_g5v0d10v5_TNBBPH_1 N4 CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5_TNBBPH
Xsky130_fd_pr__nfet_g5v0d10v5_TNBBPH_2 VSS CMFB N4 VSS sky130_fd_pr__nfet_g5v0d10v5_TNBBPH
Xsky130_fd_pr__nfet_g5v0d10v5_TNBBPH_3 VSS CMFB N3 VSS sky130_fd_pr__nfet_g5v0d10v5_TNBBPH
Xsky130_fd_pr__nfet_g5v0d10v5_TNWANH_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_TNWANH
Xsky130_fd_pr__nfet_g5v0d10v5_TNWANH_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_TNWANH
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_0 VCC out Vb2 N2 sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_2 VCC N2 Vb2 out sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_1 VCC N1 Vb2 out2 sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_3 VCC out2 Vb2 N1 sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7
Xsky130_fd_pr__nfet_g5v0d10v5_NYY6SB_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_NYY6SB
Xsky130_fd_pr__nfet_g5v0d10v5_NYY6SB_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_NYY6SB
Xsky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7
Xsky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7
Xsky130_fd_pr__pfet_g5v0d10v5_DEERZ7_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_DEERZ7
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_0 N4 Vb3 out VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0
Xsky130_fd_pr__pfet_g5v0d10v5_DEERZ7_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_DEERZ7
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_1 out2 Vb3 N3 VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_2 out Vb3 N4 VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0
Xsky130_fd_pr__pfet_g5v0d10v5_JEERZ7_0 VCC N1 Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VK4LZ7 a_n108_n836# a_n50_n862# w_n144_n898#
+ a_50_n836#
X0 a_50_n836# a_n50_n862# a_n108_n836# w_n144_n898# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0 a_n108_n50# a_50_n50# a_n50_n76# VSUBS
X0 a_50_n50# a_n50_n76# a_n108_n50# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7 a_50_n800# a_n50_n826# a_n108_n800# w_n144_n862#
X0 a_50_n800# a_n50_n826# a_n108_n800# w_n144_n862# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SAT828 a_n108_n769# a_n50_n857# a_50_n769# VSUBS
X0 a_50_n769# a_n50_n857# a_n108_n769# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GUWUK4#0 a_n108_n19# a_n50_n107# a_50_n19# VSUBS
X0 a_50_n19# a_n50_n107# a_n108_n19# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0 w_n144_n162# a_50_n100# a_n50_n126#
+ a_n108_n100#
X0 a_50_n100# a_n50_n126# a_n108_n100# w_n144_n162# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SAC338 a_50_n800# a_n50_n826# a_n108_n800# VSUBS
X0 a_50_n800# a_n50_n826# a_n108_n800# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.6 as=2.32 ps=16.6 w=8 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7#0 a_50_n136# a_n108_n136# a_n50_n162#
+ w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt input_stage Vb5 Vb1 INP N4 N3 INN N2 N1 VCC VSS
Xsky130_fd_pr__pfet_g5v0d10v5_VK4LZ7_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_VK4LZ7
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_0 VSS m1_n402_n3947# Vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_1 VSS m1_n402_n3947# Vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_2 m1_n402_n3947# VSS Vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_3 m1_n402_n3947# VSS Vb5 VSS sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0
Xsky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_1 N4 INN m1_n402_90# VCC sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7
Xsky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_0 N3 INP m1_n402_90# VCC sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7
Xsky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_2 m1_n402_90# INN N4 VCC sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7
Xsky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_3 m1_n402_90# INP N3 VCC sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7
Xsky130_fd_pr__nfet_g5v0d10v5_SAT828_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_SAT828
Xsky130_fd_pr__nfet_g5v0d10v5_GUWUK4_0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_GUWUK4#0
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_0 VCC m1_n402_90# Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0
Xsky130_fd_pr__nfet_g5v0d10v5_SAT828_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_SAT828
Xsky130_fd_pr__nfet_g5v0d10v5_GUWUK4_1 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_GUWUK4#0
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_1 VCC m1_n402_90# Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_2 VCC VCC Vb1 m1_n402_90# sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0
Xsky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_3 VCC VCC Vb1 m1_n402_90# sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0
Xsky130_fd_pr__nfet_g5v0d10v5_SAC338_0 m1_n402_n3947# INN N2 VSS sky130_fd_pr__nfet_g5v0d10v5_SAC338
Xsky130_fd_pr__nfet_g5v0d10v5_SAC338_1 N2 INN m1_n402_n3947# VSS sky130_fd_pr__nfet_g5v0d10v5_SAC338
Xsky130_fd_pr__nfet_g5v0d10v5_SAC338_2 m1_n402_n3947# INP N1 VSS sky130_fd_pr__nfet_g5v0d10v5_SAC338
Xsky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7#0
Xsky130_fd_pr__nfet_g5v0d10v5_SAC338_3 N1 INP m1_n402_n3947# VSS sky130_fd_pr__nfet_g5v0d10v5_SAC338
Xsky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7#0
Xsky130_fd_pr__pfet_g5v0d10v5_VK4LZ7_0 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5_VK4LZ7
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_8UT6AQ a_n108_n81# a_50_n81# a_n50_n107# VSUBS
X0 a_50_n81# a_n50_n107# a_n108_n81# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt total VCC VSS INP INN VOUT
Xsky130_fd_pr__nfet_g5v0d10v5_VNB5GC_1 VSS m1_6795_368# diff_to_single_ended_1/v VSS
+ sky130_fd_pr__nfet_g5v0d10v5_VNB5GC
Xcurrent_source_0 input_stage_0/Vb5 VSS folded_cascode_0/Vb3 folded_cascode_0/Vb2
+ cmfb_block_0/Vb1 VCC current_source
Xcmfb_block_0 cmfb_block_0/Vb1 cmfb_block_0/CMFB cmfb_block_0/VREF cmfb_block_0/IP
+ VCC VSS cmfb_block_0/IN cmfb_block
Xsky130_fd_pr__cap_mim_m3_1_N2QRHY_0 VSS cmfb_block_0/CMFB sky130_fd_pr__cap_mim_m3_1_N2QRHY
Xsky130_fd_pr__pfet_g5v0d10v5_2V6JZ7_0 VCC VOUT VCC m1_6795_368# sky130_fd_pr__pfet_g5v0d10v5_2V6JZ7
Xsky130_fd_pr__pfet_g5v0d10v5_GX3LZ5_0 VCC diff_to_single_ended_1/v m1_6795_368# VCC
+ sky130_fd_pr__pfet_g5v0d10v5_GX3LZ5
Xdiff_to_single_ended_1 cmfb_block_0/IN input_stage_0/Vb5 diff_to_single_ended_1/v
+ cmfb_block_0/IP VCC VSS diff_to_single_ended
Xsky130_fd_pr__nfet_g5v0d10v5_TNTUPH_0 cmfb_block_0/VREF VCC VCC VSS sky130_fd_pr__nfet_g5v0d10v5_TNTUPH#0
Xfolded_cascode_0 folded_cascode_0/Vb3 folded_cascode_0/Vb2 cmfb_block_0/Vb1 cmfb_block_0/CMFB
+ cmfb_block_0/IN input_stage_0/N4 input_stage_0/N3 input_stage_0/N2 cmfb_block_0/IP
+ input_stage_0/N1 VCC VSS folded_cascode
Xinput_stage_0 input_stage_0/Vb5 cmfb_block_0/Vb1 INP input_stage_0/N4 input_stage_0/N3
+ INN input_stage_0/N2 input_stage_0/N1 VCC VSS input_stage
Xsky130_fd_pr__nfet_g5v0d10v5_8UT6AQ_0 VSS cmfb_block_0/VREF cmfb_block_0/VREF VSS
+ sky130_fd_pr__nfet_g5v0d10v5_8UT6AQ
Xsky130_fd_pr__nfet_g5v0d10v5_NY97Z6_0 VOUT m1_6795_368# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_NY97Z6
.ends

