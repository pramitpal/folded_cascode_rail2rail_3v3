magic
tech sky130A
magscale 1 2
timestamp 1697281155
<< nwell >>
rect 2178 -1823 4555 634
<< mvpsubdiff >>
rect 2301 -1934 2349 -1910
rect 2301 -2096 2307 -1934
rect 2343 -2096 2349 -1934
rect 4383 -1934 4431 -1910
rect 2301 -2120 2349 -2096
rect 4383 -2096 4389 -1934
rect 4425 -2096 4431 -1934
rect 4383 -2120 4431 -2096
<< mvnsubdiff >>
rect 2301 460 2349 501
rect 2301 -1698 2308 460
rect 2342 -1698 2349 460
rect 4383 460 4431 501
rect 2301 -1732 2349 -1698
rect 4383 -1698 4390 460
rect 4424 -1698 4431 460
rect 4383 -1732 4431 -1698
<< mvpsubdiffcont >>
rect 2307 -2096 2343 -1934
rect 4389 -2096 4425 -1934
<< mvnsubdiffcont >>
rect 2308 -1698 2342 460
rect 4390 -1698 4424 460
<< poly >>
rect 2949 354 3049 401
rect 2949 320 2965 354
rect 3033 320 3049 354
rect 2949 304 3049 320
rect 3237 354 3337 401
rect 3237 320 3253 354
rect 3321 320 3337 354
rect 3237 304 3337 320
rect 3395 354 3495 401
rect 3395 320 3411 354
rect 3479 320 3495 354
rect 3395 304 3495 320
rect 3683 354 3783 401
rect 3683 320 3699 354
rect 3767 320 3783 354
rect 3683 304 3783 320
rect 2949 -612 3049 -565
rect 2949 -646 2965 -612
rect 3033 -646 3049 -612
rect 2949 -662 3049 -646
rect 3237 -612 3337 -565
rect 3237 -646 3253 -612
rect 3321 -646 3337 -612
rect 3237 -662 3337 -646
rect 3395 -612 3495 -565
rect 3395 -646 3411 -612
rect 3479 -646 3495 -612
rect 3395 -662 3495 -646
rect 3683 -612 3783 -565
rect 3683 -646 3699 -612
rect 3767 -646 3783 -612
rect 3683 -662 3783 -646
rect 2949 -850 3049 -834
rect 2949 -884 2965 -850
rect 3033 -884 3049 -850
rect 2949 -931 3049 -884
rect 3237 -850 3337 -834
rect 3237 -884 3253 -850
rect 3321 -884 3337 -850
rect 3237 -931 3337 -884
rect 3395 -850 3495 -834
rect 3395 -884 3411 -850
rect 3479 -884 3495 -850
rect 3395 -931 3495 -884
rect 3683 -850 3783 -834
rect 3683 -884 3699 -850
rect 3767 -884 3783 -850
rect 3683 -931 3783 -884
rect 2761 -1864 2961 -1848
rect 2761 -1898 2777 -1864
rect 2945 -1898 2961 -1864
rect 2761 -1936 2961 -1898
rect 3137 -1864 3337 -1848
rect 3137 -1898 3153 -1864
rect 3321 -1898 3337 -1864
rect 3137 -1936 3337 -1898
rect 3395 -1864 3595 -1848
rect 3395 -1898 3411 -1864
rect 3579 -1898 3595 -1864
rect 3395 -1936 3595 -1898
rect 3771 -1864 3971 -1848
rect 3771 -1898 3787 -1864
rect 3955 -1898 3971 -1864
rect 3771 -1936 3971 -1898
<< polycont >>
rect 2965 320 3033 354
rect 3253 320 3321 354
rect 3411 320 3479 354
rect 3699 320 3767 354
rect 2965 -646 3033 -612
rect 3253 -646 3321 -612
rect 3411 -646 3479 -612
rect 3699 -646 3767 -612
rect 2965 -884 3033 -850
rect 3253 -884 3321 -850
rect 3411 -884 3479 -850
rect 3699 -884 3767 -850
rect 2777 -1898 2945 -1864
rect 3153 -1898 3321 -1864
rect 3411 -1898 3579 -1864
rect 3787 -1898 3955 -1864
<< locali >>
rect 2415 548 4317 582
rect 2301 489 2349 501
rect 2415 489 2449 548
rect 2301 460 2449 489
rect 2773 469 2807 548
rect 2301 -1698 2308 460
rect 2342 413 2449 460
rect 2903 444 2937 548
rect 3349 413 3383 548
rect 3795 422 3829 548
rect 3925 476 3959 548
rect 4283 489 4317 548
rect 4383 489 4431 501
rect 4283 460 4431 489
rect 4283 413 4390 460
rect 2342 223 2349 413
rect 2415 401 2449 413
rect 4283 401 4317 413
rect 2949 320 2965 354
rect 3033 320 3253 354
rect 3321 320 3411 354
rect 3479 320 3699 354
rect 3767 320 3783 354
rect 2415 282 2807 316
rect 2415 226 2449 282
rect 2773 232 2807 282
rect 3925 282 4317 316
rect 3925 229 3959 282
rect 4283 223 4317 282
rect 4383 223 4390 413
rect 2342 -552 2420 223
rect 2342 -943 2349 -552
rect 4283 -553 4390 223
rect 2949 -646 2965 -612
rect 3033 -646 3130 -612
rect 3237 -646 3253 -612
rect 3321 -646 3411 -612
rect 3479 -646 3495 -612
rect 3596 -646 3699 -612
rect 3767 -646 3783 -612
rect 3347 -850 3381 -646
rect 2415 -884 2807 -850
rect 2949 -884 2965 -850
rect 3033 -884 3129 -850
rect 3237 -884 3253 -850
rect 3321 -884 3411 -850
rect 3479 -884 3495 -850
rect 3597 -884 3699 -850
rect 3767 -884 3783 -850
rect 3925 -884 4317 -849
rect 2415 -943 2449 -884
rect 2773 -943 2807 -884
rect 2342 -946 2449 -943
rect 2342 -1698 2441 -946
rect 3925 -960 3960 -884
rect 4282 -943 4317 -884
rect 4383 -943 4390 -553
rect 4282 -966 4390 -943
rect 2301 -1719 2441 -1698
rect 4283 -1698 4390 -966
rect 4424 -1698 4431 460
rect 2301 -1732 2349 -1719
rect 3191 -1864 3225 -1710
rect 3507 -1864 3541 -1708
rect 4283 -1719 4431 -1698
rect 4383 -1732 4431 -1719
rect 2761 -1898 2777 -1864
rect 2945 -1898 2961 -1864
rect 3137 -1898 3153 -1864
rect 3321 -1898 3337 -1864
rect 3395 -1898 3411 -1864
rect 3579 -1898 3595 -1864
rect 3771 -1898 3787 -1864
rect 3955 -1898 3971 -1864
rect 2301 -1934 2349 -1910
rect 2301 -2096 2307 -1934
rect 2343 -1948 2349 -1934
rect 4383 -1934 4431 -1910
rect 4383 -1948 4389 -1934
rect 2343 -2014 2458 -1948
rect 2343 -2024 2473 -2014
rect 2343 -2096 2349 -2024
rect 2301 -2120 2349 -2096
rect 2439 -2074 2473 -2024
rect 2597 -2074 2631 -1959
rect 2972 -2074 3006 -1997
rect 3349 -2074 3383 -1998
rect 3726 -2074 3760 -1978
rect 4101 -2074 4135 -2020
rect 4259 -2024 4389 -1948
rect 4259 -2074 4293 -2024
rect 2439 -2108 4293 -2074
rect 4383 -2096 4389 -2024
rect 4425 -2096 4431 -1934
rect 4383 -2120 4431 -2096
<< viali >>
rect 3130 -646 3164 -612
rect 3562 -646 3596 -612
rect 3129 -884 3163 -850
rect 3563 -884 3597 -850
rect 2777 -1898 2945 -1864
rect 3787 -1898 3955 -1864
<< metal1 >>
rect 3061 194 3095 435
rect 3191 416 3225 443
rect 3507 416 3541 443
rect 3182 410 3234 416
rect 3182 352 3234 358
rect 3498 410 3550 416
rect 3498 352 3550 358
rect 3637 198 3671 441
rect 2903 -1661 2937 -481
rect 3061 -689 3095 -494
rect 3191 -509 3225 -506
rect 3182 -515 3234 -509
rect 3182 -573 3234 -567
rect 3124 -612 3170 -600
rect 3250 -612 3256 -603
rect 3124 -646 3130 -612
rect 3164 -646 3256 -612
rect 3124 -658 3170 -646
rect 3250 -655 3256 -646
rect 3308 -655 3314 -603
rect 3349 -689 3383 -449
rect 3507 -515 3541 -486
rect 3492 -567 3498 -515
rect 3550 -567 3556 -515
rect 3421 -603 3473 -597
rect 3550 -612 3608 -606
rect 3473 -646 3562 -612
rect 3596 -646 3608 -612
rect 3550 -652 3608 -646
rect 3421 -661 3473 -655
rect 3636 -689 3670 -518
rect 3061 -723 3670 -689
rect 3052 -758 3104 -752
rect 3628 -758 3680 -752
rect 3104 -801 3628 -767
rect 3052 -816 3104 -810
rect 3061 -964 3095 -816
rect 3123 -850 3169 -838
rect 3256 -850 3262 -841
rect 3123 -884 3129 -850
rect 3163 -884 3262 -850
rect 3123 -896 3169 -884
rect 3256 -893 3262 -884
rect 3314 -893 3320 -841
rect 3176 -983 3182 -931
rect 3234 -983 3240 -931
rect 3191 -992 3225 -983
rect 2903 -1719 2938 -1661
rect 3191 -1679 3225 -1609
rect 2904 -1854 2938 -1719
rect 3176 -1731 3182 -1679
rect 3234 -1731 3240 -1679
rect 3349 -1719 3383 -801
rect 3628 -816 3680 -810
rect 3414 -841 3466 -835
rect 3551 -850 3609 -844
rect 3466 -884 3563 -850
rect 3597 -884 3609 -850
rect 3551 -890 3609 -884
rect 3414 -899 3466 -893
rect 3498 -931 3550 -925
rect 3498 -989 3550 -983
rect 3507 -993 3541 -989
rect 3637 -1004 3671 -816
rect 3507 -1679 3541 -1662
rect 3492 -1731 3498 -1679
rect 3550 -1731 3556 -1679
rect 2715 -1864 2957 -1854
rect 3795 -1855 3829 -419
rect 3775 -1864 3964 -1855
rect 2715 -1898 2777 -1864
rect 2945 -1898 3787 -1864
rect 3955 -1898 4017 -1864
rect 2715 -1908 2957 -1898
rect 3775 -1908 4017 -1898
rect 2715 -2024 2749 -1908
rect 3077 -1988 3083 -1936
rect 3135 -1988 3141 -1936
rect 3592 -1988 3598 -1936
rect 3650 -1988 3656 -1936
rect 3983 -1961 4017 -1908
rect 3092 -2004 3126 -1988
rect 3091 -2075 3125 -2015
rect 3607 -2075 3641 -1988
rect 3091 -2109 3641 -2075
<< via1 >>
rect 3182 358 3234 410
rect 3498 358 3550 410
rect 3182 -567 3234 -515
rect 3256 -655 3308 -603
rect 3498 -567 3550 -515
rect 3421 -655 3473 -603
rect 3052 -810 3104 -758
rect 3262 -893 3314 -841
rect 3182 -983 3234 -931
rect 3182 -1731 3234 -1679
rect 3628 -810 3680 -758
rect 3414 -893 3466 -841
rect 3498 -983 3550 -931
rect 3498 -1731 3550 -1679
rect 3083 -1988 3135 -1936
rect 3598 -1988 3650 -1936
<< metal2 >>
rect 3178 414 3238 423
rect 3494 414 3554 423
rect 3176 358 3178 410
rect 3238 358 3240 410
rect 3492 358 3494 410
rect 3554 358 3556 410
rect 3178 345 3238 354
rect 3494 345 3554 354
rect 3498 -515 3550 -509
rect 3176 -567 3182 -515
rect 3234 -567 3240 -515
rect 2767 -601 2823 -592
rect 2218 -646 2767 -612
rect 2767 -666 2823 -657
rect 3048 -754 3108 -745
rect 3046 -810 3048 -758
rect 3108 -810 3110 -758
rect 3048 -823 3108 -814
rect 2766 -839 2822 -830
rect 2218 -884 2766 -850
rect 2766 -904 2822 -895
rect 3191 -925 3225 -567
rect 3498 -573 3550 -567
rect 3256 -599 3479 -597
rect 3256 -603 3337 -599
rect 3308 -655 3337 -603
rect 3256 -659 3337 -655
rect 3397 -603 3479 -599
rect 3397 -655 3421 -603
rect 3473 -655 3479 -603
rect 3397 -659 3479 -655
rect 3256 -661 3479 -659
rect 3262 -837 3472 -835
rect 3262 -841 3336 -837
rect 3314 -893 3336 -841
rect 3262 -897 3336 -893
rect 3396 -841 3472 -837
rect 3396 -893 3414 -841
rect 3466 -893 3472 -841
rect 3396 -897 3472 -893
rect 3262 -899 3472 -897
rect 3182 -931 3234 -925
rect 3507 -931 3541 -573
rect 3624 -754 3684 -745
rect 3622 -810 3624 -758
rect 3684 -810 3686 -758
rect 3624 -823 3684 -814
rect 3492 -983 3498 -931
rect 3550 -983 3556 -931
rect 3182 -989 3234 -983
rect 3182 -1679 3234 -1673
rect 3092 -1722 3182 -1688
rect 3092 -1930 3126 -1722
rect 3182 -1737 3234 -1731
rect 3498 -1679 3550 -1673
rect 3550 -1722 3641 -1688
rect 3498 -1737 3550 -1731
rect 3607 -1930 3641 -1722
rect 3083 -1936 3135 -1930
rect 3083 -1994 3135 -1988
rect 3598 -1936 3650 -1930
rect 3598 -1994 3650 -1988
<< via2 >>
rect 3178 410 3238 414
rect 3494 410 3554 414
rect 3178 358 3182 410
rect 3182 358 3234 410
rect 3234 358 3238 410
rect 3494 358 3498 410
rect 3498 358 3550 410
rect 3550 358 3554 410
rect 3178 354 3238 358
rect 3494 354 3554 358
rect 2767 -657 2823 -601
rect 3048 -758 3108 -754
rect 3048 -810 3052 -758
rect 3052 -810 3104 -758
rect 3104 -810 3108 -758
rect 3048 -814 3108 -810
rect 2766 -895 2822 -839
rect 3337 -659 3397 -599
rect 3336 -897 3396 -837
rect 3624 -758 3684 -754
rect 3624 -810 3628 -758
rect 3628 -810 3680 -758
rect 3680 -810 3684 -758
rect 3624 -814 3684 -810
<< metal3 >>
rect 3173 414 3243 419
rect 3173 354 3178 414
rect 3238 354 3243 414
rect 3173 349 3243 354
rect 3489 414 3559 419
rect 3489 354 3494 414
rect 3554 354 3559 414
rect 3489 349 3559 354
rect 3178 -311 3238 349
rect 3048 -371 3238 -311
rect 3494 -311 3554 349
rect 3494 -371 3684 -311
rect 2762 -599 2828 -596
rect 2894 -597 2958 -591
rect 2762 -601 2894 -599
rect 2762 -657 2767 -601
rect 2823 -657 2894 -601
rect 2762 -659 2894 -657
rect 2762 -662 2828 -659
rect 2894 -667 2958 -661
rect 3048 -749 3108 -371
rect 3191 -661 3197 -597
rect 3261 -599 3267 -597
rect 3332 -599 3402 -594
rect 3261 -659 3337 -599
rect 3397 -659 3402 -599
rect 3261 -661 3267 -659
rect 3332 -664 3402 -659
rect 3624 -749 3684 -371
rect 3043 -754 3113 -749
rect 3043 -814 3048 -754
rect 3108 -814 3113 -754
rect 3043 -819 3113 -814
rect 3619 -754 3689 -749
rect 3619 -814 3624 -754
rect 3684 -814 3689 -754
rect 3619 -819 3689 -814
rect 2761 -837 2827 -834
rect 2894 -835 2958 -829
rect 2761 -839 2894 -837
rect 2761 -895 2766 -839
rect 2822 -895 2894 -839
rect 2761 -897 2894 -895
rect 2761 -900 2827 -897
rect 3191 -899 3197 -835
rect 3261 -837 3267 -835
rect 3331 -837 3401 -832
rect 3261 -897 3336 -837
rect 3396 -897 3401 -837
rect 3261 -899 3267 -897
rect 2894 -905 2958 -899
rect 3331 -902 3401 -897
<< via3 >>
rect 2894 -661 2958 -597
rect 3197 -661 3261 -597
rect 2894 -899 2958 -835
rect 3197 -899 3261 -835
<< metal4 >>
rect 2893 -597 2959 -596
rect 2893 -661 2894 -597
rect 2958 -599 2959 -597
rect 3196 -597 3262 -596
rect 3196 -599 3197 -597
rect 2958 -659 3197 -599
rect 2958 -661 2959 -659
rect 2893 -662 2959 -661
rect 3196 -661 3197 -659
rect 3261 -661 3262 -597
rect 3196 -662 3262 -661
rect 2893 -835 2959 -834
rect 2893 -899 2894 -835
rect 2958 -837 2959 -835
rect 3196 -835 3262 -834
rect 3196 -837 3197 -835
rect 2958 -897 3197 -837
rect 2958 -899 2959 -897
rect 2893 -900 2959 -899
rect 3196 -899 3197 -897
rect 3261 -899 3262 -835
rect 3196 -900 3262 -899
use sky130_fd_pr__nfet_g5v0d10v5_6DL6AA  sky130_fd_pr__nfet_g5v0d10v5_6DL6AA_0
timestamp 1697281155
transform 1 0 3237 0 1 -1986
box -158 -76 158 76
use sky130_fd_pr__nfet_g5v0d10v5_6DL6AA  sky130_fd_pr__nfet_g5v0d10v5_6DL6AA_1
timestamp 1697281155
transform 1 0 2861 0 1 -1986
box -158 -76 158 76
use sky130_fd_pr__nfet_g5v0d10v5_6DL6AA  sky130_fd_pr__nfet_g5v0d10v5_6DL6AA_2
timestamp 1697281155
transform 1 0 3495 0 1 -1986
box -158 -76 158 76
use sky130_fd_pr__nfet_g5v0d10v5_6DL6AA  sky130_fd_pr__nfet_g5v0d10v5_6DL6AA_3
timestamp 1697281155
transform 1 0 3871 0 1 -1986
box -158 -76 158 76
use sky130_fd_pr__nfet_g5v0d10v5_GUWUK4  sky130_fd_pr__nfet_g5v0d10v5_GUWUK4_0
timestamp 1697281155
transform 1 0 2535 0 1 -2017
box -108 -107 108 107
use sky130_fd_pr__nfet_g5v0d10v5_GUWUK4  sky130_fd_pr__nfet_g5v0d10v5_GUWUK4_1
timestamp 1697281155
transform 1 0 4197 0 1 -2017
box -108 -107 108 107
use sky130_fd_pr__pfet_g5v0d10v5_3JERZF  sky130_fd_pr__pfet_g5v0d10v5_3JERZF_0
timestamp 1697281155
transform 1 0 2611 0 1 -1295
box -274 -502 274 464
use sky130_fd_pr__pfet_g5v0d10v5_3JERZF  sky130_fd_pr__pfet_g5v0d10v5_3JERZF_1
timestamp 1697281155
transform 1 0 4121 0 1 -1295
box -274 -502 274 464
use sky130_fd_pr__pfet_g5v0d10v5_3JERZF  sky130_fd_pr__pfet_g5v0d10v5_3JERZF_2
timestamp 1697281155
transform 1 0 2611 0 1 -129
box -274 -502 274 464
use sky130_fd_pr__pfet_g5v0d10v5_3JERZF  sky130_fd_pr__pfet_g5v0d10v5_3JERZF_3
timestamp 1697281155
transform 1 0 4121 0 1 -129
box -274 -502 274 464
use sky130_fd_pr__pfet_g5v0d10v5_6LM9S7  sky130_fd_pr__pfet_g5v0d10v5_6LM9S7_4
timestamp 1697281155
transform 1 0 3733 0 1 451
box -174 -116 174 116
use sky130_fd_pr__pfet_g5v0d10v5_6LM9S7  sky130_fd_pr__pfet_g5v0d10v5_6LM9S7_5
timestamp 1697281155
transform 1 0 3445 0 1 451
box -174 -116 174 116
use sky130_fd_pr__pfet_g5v0d10v5_6LM9S7  sky130_fd_pr__pfet_g5v0d10v5_6LM9S7_6
timestamp 1697281155
transform 1 0 3287 0 1 451
box -174 -116 174 116
use sky130_fd_pr__pfet_g5v0d10v5_6LM9S7  sky130_fd_pr__pfet_g5v0d10v5_6LM9S7_7
timestamp 1697281155
transform 1 0 2999 0 1 451
box -174 -116 174 116
use sky130_fd_pr__pfet_g5v0d10v5_7JP9SF  sky130_fd_pr__pfet_g5v0d10v5_7JP9SF_0
timestamp 1697281155
transform 1 0 2611 0 1 487
box -274 -152 274 114
use sky130_fd_pr__pfet_g5v0d10v5_7JP9SF  sky130_fd_pr__pfet_g5v0d10v5_7JP9SF_1
timestamp 1697281155
transform 1 0 4121 0 1 487
box -274 -152 274 114
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_8
timestamp 1697281155
transform 1 0 3733 0 1 -1331
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_9
timestamp 1697281155
transform 1 0 2999 0 1 -1331
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_10
timestamp 1697281155
transform 1 0 3287 0 1 -1331
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_11
timestamp 1697281155
transform 1 0 3445 0 1 -1331
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_12
timestamp 1697281155
transform 1 0 3733 0 1 -165
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_13
timestamp 1697281155
transform 1 0 2999 0 1 -165
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_14
timestamp 1697281155
transform 1 0 3287 0 1 -165
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_15
timestamp 1697281155
transform 1 0 3445 0 1 -165
box -174 -466 174 466
<< labels >>
flabel locali s 3602 329 3602 329 0 FreeSans 800 0 0 0 Vb1
flabel locali s 3614 -633 3614 -633 0 FreeSans 800 0 0 0 IN
flabel locali s 3620 -861 3620 -861 0 FreeSans 800 0 0 0 IP
flabel locali s 3446 568 3446 568 0 FreeSans 800 0 0 0 VCC
flabel locali s 2680 -2095 2680 -2095 0 FreeSans 800 0 0 0 VSS
flabel metal2 s 3622 -1846 3622 -1846 0 FreeSans 800 0 0 0 CMFB
flabel locali s 3364 -744 3364 -744 0 FreeSans 800 0 0 0 VREF
<< end >>
