magic
tech sky130A
timestamp 1697284980
<< error_p >>
rect -87 431 87 433
rect -87 -431 -72 431
rect -54 398 54 400
rect -54 -398 -39 398
rect 39 -398 54 398
rect -54 -400 54 -398
rect 72 -431 87 431
rect -87 -433 87 -431
<< nwell >>
rect -72 -431 72 431
<< mvpmos >>
rect -25 -400 25 400
<< mvpdiff >>
rect -54 394 -25 400
rect -54 -394 -48 394
rect -31 -394 -25 394
rect -54 -400 -25 -394
rect 25 394 54 400
rect 25 -394 31 394
rect 48 -394 54 394
rect 25 -400 54 -394
<< mvpdiffc >>
rect -48 -394 -31 394
rect 31 -394 48 394
<< poly >>
rect -25 400 25 413
rect -25 -413 25 -400
<< locali >>
rect -48 394 -31 402
rect -48 -402 -31 -394
rect 31 394 48 402
rect 31 -402 48 -394
<< viali >>
rect -48 -394 -31 394
rect 31 -394 48 394
<< metal1 >>
rect -51 394 -28 400
rect -51 -394 -48 394
rect -31 -394 -28 394
rect -51 -400 -28 -394
rect 28 394 51 400
rect 28 -394 31 394
rect 48 -394 51 394
rect 28 -400 51 -394
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
