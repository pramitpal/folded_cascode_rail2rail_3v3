magic
tech sky130A
magscale 1 2
timestamp 1698929273
<< nwell >>
rect -656 2791 6236 4738
<< mvpsubdiff >>
rect -582 2610 -534 2654
rect -582 48 -576 2610
rect -540 48 -534 2610
rect -582 14 -534 48
rect 4764 2600 4812 2644
rect 4764 38 4770 2600
rect 4806 38 4812 2600
rect 4764 4 4812 38
rect 6122 2600 6170 2644
rect 6122 38 6128 2600
rect 6164 38 6170 2600
rect 6122 4 6170 38
<< mvnsubdiff >>
rect 4776 4566 4824 4596
rect -582 4530 -534 4560
rect -582 2996 -576 4530
rect -540 2996 -534 4530
rect -582 2926 -534 2996
rect 4776 3032 4782 4566
rect 4818 3032 4824 4566
rect 4776 2962 4824 3032
rect 6122 4566 6170 4596
rect 6122 3032 6128 4566
rect 6164 3032 6170 4566
rect 6122 2962 6170 3032
<< mvpsubdiffcont >>
rect -576 48 -540 2610
rect 4770 38 4806 2600
rect 6128 38 6164 2600
<< mvnsubdiffcont >>
rect -576 2996 -540 4530
rect 4782 3032 4818 4566
rect 6128 3032 6164 4566
<< poly >>
rect -378 3739 22 3786
rect -378 3705 -362 3739
rect 6 3705 22 3739
rect -378 3689 22 3705
rect 210 3739 610 3786
rect 210 3705 226 3739
rect 594 3705 610 3739
rect 210 3689 610 3705
rect 798 3739 1198 3786
rect 798 3705 814 3739
rect 1182 3705 1198 3739
rect 798 3689 1198 3705
rect 1386 3739 1786 3786
rect 1386 3705 1402 3739
rect 1770 3705 1786 3739
rect 1386 3689 1786 3705
rect 1974 3739 2374 3786
rect 1974 3705 1990 3739
rect 2358 3705 2374 3739
rect 1974 3689 2374 3705
rect 2432 3739 2832 3786
rect 2432 3705 2448 3739
rect 2816 3705 2832 3739
rect 2432 3689 2832 3705
rect 3020 3739 3420 3786
rect 3020 3705 3036 3739
rect 3404 3705 3420 3739
rect 3020 3689 3420 3705
rect 3608 3739 4008 3786
rect 3608 3705 3624 3739
rect 3992 3705 4008 3739
rect 3608 3689 4008 3705
rect 4196 3739 4596 3786
rect 4196 3705 4212 3739
rect 4580 3705 4596 3739
rect 4196 3689 4596 3705
<< polycont >>
rect -362 3705 6 3739
rect 226 3705 594 3739
rect 814 3705 1182 3739
rect 1402 3705 1770 3739
rect 1990 3705 2358 3739
rect 2448 3705 2816 3739
rect 3036 3705 3404 3739
rect 3624 3705 3992 3739
rect 4212 3705 4580 3739
<< locali >>
rect 4776 4568 4824 4596
rect 4620 4566 4972 4568
rect -582 4532 -534 4560
rect -582 4530 -410 4532
rect -582 2996 -576 4530
rect -540 3850 -410 4530
rect -540 3739 -390 3850
rect 34 3739 68 3818
rect -540 3705 -362 3739
rect 6 3705 68 3739
rect 164 3739 198 3850
rect 622 3739 656 3818
rect 1928 3739 1962 3793
rect 2844 3739 2878 3847
rect 4150 3739 4184 3802
rect 4620 3797 4782 4566
rect 4608 3739 4782 3797
rect 164 3705 226 3739
rect 594 3705 656 3739
rect 798 3705 814 3739
rect 1182 3705 1402 3739
rect 1770 3705 1990 3739
rect 2358 3705 2448 3739
rect 2816 3705 3036 3739
rect 3404 3705 3624 3739
rect 3992 3705 4008 3739
rect 4150 3705 4212 3739
rect 4580 3705 4782 3739
rect -540 2996 -390 3705
rect 622 3501 656 3705
rect 2386 3521 2420 3705
rect 4608 3433 4782 3705
rect 4620 3038 4782 3433
rect -582 2926 -534 2996
rect -424 2923 -390 2996
rect 34 2923 68 3031
rect 1928 2923 1962 2985
rect 2844 2923 2878 3027
rect 4150 2923 4184 3037
rect 4608 2923 4642 3037
rect 4776 3032 4782 3038
rect 4818 3038 4972 4566
rect 4818 3032 4824 3038
rect 4776 2962 4824 3032
rect -424 2889 68 2923
rect 226 2728 595 2922
rect 1085 2889 3696 2923
rect 4150 2889 4642 2923
rect 4951 2939 4985 3014
rect 5397 3000 5559 4574
rect 6122 4566 6170 4596
rect 6122 4546 6128 4566
rect 5109 2939 5143 2993
rect 4951 2905 5143 2939
rect 5239 2939 5273 3000
rect 5397 2998 5561 3000
rect 5527 2939 5561 2998
rect 5815 2939 5849 3041
rect 5980 3032 6128 4546
rect 6164 3032 6170 4566
rect 5980 3030 6170 3032
rect 5973 2939 6007 2996
rect 6122 2962 6170 3030
rect 5239 2905 5347 2939
rect 5527 2905 5617 2939
rect 5815 2905 6007 2939
rect 2386 2824 2420 2889
rect 1792 2810 1838 2816
rect 1792 2776 1795 2810
rect 1835 2776 1838 2810
rect 2968 2810 3014 2816
rect 1792 2728 1838 2776
rect 2968 2776 2971 2810
rect 3011 2776 3014 2810
rect 2968 2728 3014 2776
rect 5239 2728 5273 2787
rect -424 2694 68 2728
rect 226 2694 3687 2728
rect 4150 2694 4642 2728
rect -582 2610 -534 2654
rect -424 2612 -390 2694
rect -582 48 -576 2610
rect -540 2604 -534 2610
rect -540 1675 -412 2604
rect 34 1856 68 2694
rect 1798 2614 1832 2694
rect 2974 2620 3008 2694
rect 164 1675 198 1896
rect 1340 1675 1374 1908
rect 3432 1675 3466 1890
rect 4150 1874 4184 2694
rect 4608 2631 4642 2694
rect 4951 2681 5143 2715
rect 4764 2631 4812 2644
rect 4951 2631 4985 2681
rect 4608 2630 4985 2631
rect 4608 2600 4968 2630
rect 5109 2623 5143 2681
rect 5239 2694 5319 2728
rect 5239 2623 5273 2694
rect 5527 2681 5719 2715
rect 4608 2597 4770 2600
rect 4618 1675 4770 2597
rect -540 1641 68 1675
rect 164 1641 350 1675
rect 805 1641 4008 1675
rect 4150 1641 4770 1675
rect -540 1561 -390 1641
rect 34 1580 68 1641
rect 1340 1599 1374 1641
rect 3432 1579 3466 1641
rect -540 48 -412 1561
rect 4150 1553 4184 1641
rect 4608 1557 4770 1641
rect 1035 438 1081 444
rect 1035 404 1038 438
rect 1078 404 1081 438
rect -582 14 -534 48
rect 901 -40 935 90
rect 1035 74 1081 404
rect 1632 438 1678 444
rect 1632 404 1635 438
rect 1675 404 1678 438
rect 1496 -40 1530 88
rect 1632 72 1678 404
rect 3130 438 3176 444
rect 3130 404 3133 438
rect 3173 404 3176 438
rect 3130 75 3176 404
rect 3724 438 3770 444
rect 3724 404 3727 438
rect 3767 404 3770 438
rect 3282 -40 3316 88
rect 3724 66 3770 404
rect 3875 -40 3909 85
rect 4618 38 4770 1557
rect 4806 38 4968 2600
rect 5527 2583 5561 2681
rect 5685 2614 5719 2681
rect 5815 2681 6007 2715
rect 5815 2607 5849 2681
rect 5973 2620 6007 2681
rect 6122 2620 6170 2644
rect 5973 2600 6170 2620
rect 5397 2156 5431 2326
rect 5341 2122 5431 2156
rect 5397 2058 5431 2122
rect 5239 1155 5273 1328
rect 5239 1121 5431 1155
rect 5239 1061 5273 1121
rect 5397 1061 5431 1121
rect 4618 34 4968 38
rect 5973 38 6128 2600
rect 6164 38 6170 2600
rect 4764 4 4812 34
rect 5973 15 6170 38
rect 6122 4 6170 15
<< viali >>
rect -362 3705 6 3739
rect 979 3739 1013 3742
rect 226 3705 594 3739
rect 979 3705 1013 3739
rect 1402 3705 1770 3739
rect 1990 3705 2358 3739
rect 2448 3705 2816 3739
rect 3036 3705 3404 3739
rect 4212 3705 4580 3739
rect 979 3702 1013 3705
rect 1795 2776 1835 2810
rect 2386 2790 2420 2824
rect 2971 2776 3011 2810
rect 5239 2787 5273 2821
rect 1038 404 1078 438
rect 1635 404 1675 438
rect 901 -74 935 -40
rect 3133 404 3173 438
rect 3727 404 3767 438
rect 1496 -74 1530 -40
rect 3282 -74 3316 -40
rect 3875 -74 3909 -40
<< metal1 >>
rect 34 4657 6007 4691
rect 34 4538 68 4657
rect 622 4538 656 4657
rect 1210 4509 1244 4657
rect 1798 4521 1832 4657
rect 737 3994 743 4046
rect 795 3994 801 4046
rect 746 3867 792 3994
rect 1340 3878 1374 3931
rect -374 3739 18 3745
rect -374 3705 -362 3739
rect 6 3705 18 3739
rect -374 3699 18 3705
rect 214 3739 606 3745
rect 214 3705 226 3739
rect 594 3705 606 3739
rect 214 3699 606 3705
rect 161 3043 206 3100
rect 151 2991 157 3043
rect 209 2991 215 3043
rect 752 2982 786 3867
rect 1325 3826 1331 3878
rect 1383 3826 1389 3878
rect 2386 3798 2420 4657
rect 2974 4521 3008 4657
rect 3562 4542 3596 4657
rect 4150 4492 4184 4657
rect 4951 4510 4985 4657
rect 5685 4556 5719 4657
rect 5973 4531 6007 4657
rect 4005 3994 4011 4046
rect 4063 3994 4069 4046
rect 4014 3940 4060 3994
rect 3432 3878 3466 3931
rect 3417 3826 3423 3878
rect 3475 3826 3481 3878
rect 967 3748 1019 3754
rect 1019 3696 1025 3748
rect 1390 3739 1782 3745
rect 1390 3705 1402 3739
rect 1770 3705 1782 3739
rect 1390 3699 1782 3705
rect 1978 3739 2370 3745
rect 1978 3705 1990 3739
rect 2358 3705 2370 3739
rect 1978 3699 2370 3705
rect 2436 3739 2828 3745
rect 2436 3705 2448 3739
rect 2816 3705 2828 3739
rect 2436 3699 2828 3705
rect 3024 3739 3416 3745
rect 3024 3705 3036 3739
rect 3404 3705 3416 3739
rect 3024 3699 3416 3705
rect 967 3690 1019 3696
rect 1331 3663 1383 3669
rect 1331 3605 1383 3611
rect 3423 3663 3475 3669
rect 3423 3605 3475 3611
rect 1195 3141 1201 3193
rect 1253 3141 1259 3193
rect 1204 3005 1250 3141
rect 1210 2982 1244 3005
rect 1340 2982 1374 3605
rect 3432 3570 3466 3605
rect 1792 3130 1838 3244
rect 2968 3233 3014 3244
rect 3547 3141 3553 3193
rect 3605 3141 3611 3193
rect 1798 3032 1832 3130
rect 2974 3038 3008 3064
rect 3556 3044 3602 3141
rect 2965 3032 3017 3038
rect 1789 3026 1841 3032
rect 4020 2982 4054 3826
rect 4200 3739 4592 3745
rect 4200 3705 4212 3739
rect 4580 3705 4592 3739
rect 4200 3699 4592 3705
rect 2965 2974 3017 2980
rect 1789 2968 1841 2974
rect 5218 2948 5270 2954
rect 5270 2899 5311 2945
rect 5218 2890 5270 2896
rect 2377 2833 2429 2839
rect 1783 2770 1789 2822
rect 1841 2770 1847 2822
rect 2374 2784 2377 2830
rect 5233 2830 5279 2833
rect 2429 2784 2432 2830
rect 2377 2775 2429 2781
rect 2959 2770 2965 2822
rect 3017 2770 3023 2822
rect 5224 2778 5230 2830
rect 5282 2778 5288 2830
rect 5233 2775 5279 2778
rect 1789 2764 1841 2770
rect 2965 2764 3017 2770
rect 156 2645 208 2651
rect 156 2587 208 2593
rect 2371 2566 2377 2618
rect 2429 2566 2435 2618
rect 2386 2520 2420 2566
rect 1210 2304 1244 2315
rect 1195 2252 1201 2304
rect 1253 2252 1259 2304
rect 3547 2252 3553 2304
rect 3605 2252 3611 2304
rect 3426 2177 3472 2213
rect 3556 2149 3602 2252
rect 1928 2122 1962 2136
rect 1913 2070 1919 2122
rect 1971 2070 1977 2122
rect 2829 2070 2835 2122
rect 2887 2070 2893 2122
rect 1928 2050 1962 2070
rect 622 1972 656 2031
rect 2838 2029 2884 2070
rect 607 1920 613 1972
rect 665 1920 671 1972
rect 752 1925 786 1926
rect 743 1919 795 1925
rect 4020 1917 4054 1918
rect 743 1861 795 1867
rect 4011 1911 4063 1917
rect 4011 1853 4063 1859
rect 607 1534 613 1586
rect 665 1534 671 1586
rect 737 1534 743 1586
rect 795 1534 801 1586
rect 622 1499 656 1534
rect 746 1477 792 1534
rect 2371 1509 2377 1561
rect 2429 1509 2435 1561
rect 4005 1536 4011 1588
rect 4063 1536 4069 1588
rect 149 1415 155 1467
rect 207 1415 213 1467
rect 2380 1448 2426 1509
rect 4014 1477 4060 1536
rect 164 1333 198 1415
rect 622 681 656 850
rect 164 635 656 681
rect 164 585 198 635
rect 34 -40 68 49
rect 622 -40 656 635
rect 1026 398 1032 450
rect 1084 398 1090 450
rect 1032 392 1084 398
rect 895 -40 941 -28
rect 1210 -40 1244 853
rect 1623 398 1629 450
rect 1681 398 1687 450
rect 1629 392 1681 398
rect 1490 -40 1536 -28
rect 1798 -40 1832 840
rect 1928 450 1962 471
rect 1913 398 1919 450
rect 1971 398 1977 450
rect 2829 398 2835 450
rect 2887 398 2893 450
rect 1928 380 1962 398
rect 2838 341 2884 398
rect 2974 -40 3008 844
rect 3121 398 3127 450
rect 3179 398 3185 450
rect 3127 392 3179 398
rect 3276 -40 3322 -28
rect 3562 -40 3596 889
rect 3715 398 3721 450
rect 3773 398 3779 450
rect 3721 392 3773 398
rect 3869 -40 3915 -28
rect 4150 -40 4184 33
rect 4951 -40 4985 15
rect 5239 -40 5273 26
rect 5685 -40 5719 31
rect 5973 -40 6007 62
rect 34 -74 901 -40
rect 935 -74 1496 -40
rect 1530 -74 3282 -40
rect 3316 -74 3875 -40
rect 3909 -74 6007 -40
rect 895 -86 941 -74
rect 1490 -86 1536 -74
rect 3276 -86 3322 -74
rect 3869 -86 3915 -74
<< via1 >>
rect 743 3994 795 4046
rect 157 2991 209 3043
rect 1331 3826 1383 3878
rect 4011 3994 4063 4046
rect 3423 3826 3475 3878
rect 967 3742 1019 3748
rect 967 3702 979 3742
rect 979 3702 1013 3742
rect 1013 3702 1019 3742
rect 967 3696 1019 3702
rect 1331 3611 1383 3663
rect 3423 3611 3475 3663
rect 1201 3141 1253 3193
rect 3553 3141 3605 3193
rect 1789 2974 1841 3026
rect 2965 2980 3017 3032
rect 5218 2896 5270 2948
rect 1789 2810 1841 2822
rect 1789 2776 1795 2810
rect 1795 2776 1835 2810
rect 1835 2776 1841 2810
rect 1789 2770 1841 2776
rect 2377 2824 2429 2833
rect 2377 2790 2386 2824
rect 2386 2790 2420 2824
rect 2420 2790 2429 2824
rect 2377 2781 2429 2790
rect 2965 2810 3017 2822
rect 2965 2776 2971 2810
rect 2971 2776 3011 2810
rect 3011 2776 3017 2810
rect 2965 2770 3017 2776
rect 5230 2821 5282 2830
rect 5230 2787 5239 2821
rect 5239 2787 5273 2821
rect 5273 2787 5282 2821
rect 5230 2778 5282 2787
rect 156 2593 208 2645
rect 2377 2566 2429 2618
rect 1201 2252 1253 2304
rect 3553 2252 3605 2304
rect 1919 2070 1971 2122
rect 2835 2070 2887 2122
rect 613 1920 665 1972
rect 743 1867 795 1919
rect 4011 1859 4063 1911
rect 613 1534 665 1586
rect 743 1534 795 1586
rect 2377 1509 2429 1561
rect 4011 1536 4063 1588
rect 155 1415 207 1467
rect 1032 438 1084 450
rect 1032 404 1038 438
rect 1038 404 1078 438
rect 1078 404 1084 438
rect 1032 398 1084 404
rect 1629 438 1681 450
rect 1629 404 1635 438
rect 1635 404 1675 438
rect 1675 404 1681 438
rect 1629 398 1681 404
rect 1919 398 1971 450
rect 2835 398 2887 450
rect 3127 438 3179 450
rect 3127 404 3133 438
rect 3133 404 3173 438
rect 3173 404 3179 438
rect 3127 398 3179 404
rect 3721 438 3773 450
rect 3721 404 3727 438
rect 3727 404 3767 438
rect 3767 404 3773 438
rect 3721 398 3773 404
<< metal2 >>
rect 743 4046 795 4052
rect 4011 4046 4063 4052
rect 795 3997 4011 4043
rect 743 3988 795 3994
rect 4011 3988 4063 3994
rect 1331 3878 1383 3884
rect 3423 3878 3475 3884
rect 1383 3835 3423 3869
rect 1331 3820 1383 3826
rect 3423 3820 3475 3826
rect 961 3739 967 3748
rect 538 3705 967 3739
rect 157 3043 209 3049
rect 157 2985 209 2991
rect 160 2645 205 2985
rect 150 2593 156 2645
rect 208 2593 214 2645
rect 155 1467 207 1473
rect 538 1458 572 3705
rect 961 3696 967 3705
rect 1019 3696 1025 3748
rect 1340 3663 1374 3820
rect 3432 3663 3466 3820
rect 1325 3611 1331 3663
rect 1383 3611 1389 3663
rect 3417 3611 3423 3663
rect 3475 3611 3481 3663
rect 2380 3330 4113 3376
rect 1201 3193 1253 3199
rect 2380 3190 2426 3330
rect 3553 3193 3605 3199
rect 1253 3144 3553 3190
rect 1201 3135 1253 3141
rect 3553 3135 3605 3141
rect 1783 2974 1789 3026
rect 1841 2974 1847 3026
rect 2959 2980 2965 3032
rect 3017 2980 3023 3032
rect 1792 2828 1838 2974
rect 1789 2822 1841 2828
rect 2371 2781 2377 2833
rect 2429 2781 2435 2833
rect 2968 2828 3014 2980
rect 4067 2834 4113 3330
rect 5212 2945 5218 2948
rect 4444 2899 5218 2945
rect 2965 2822 3017 2828
rect 1789 2764 1841 2770
rect 2386 2624 2420 2781
rect 4051 2774 4060 2834
rect 4120 2774 4129 2834
rect 2965 2764 3017 2770
rect 2377 2618 2429 2624
rect 2377 2560 2429 2566
rect 4444 2476 4490 2899
rect 5212 2896 5218 2899
rect 5270 2896 5276 2948
rect 4626 2774 4635 2834
rect 4695 2821 4704 2834
rect 5230 2830 5282 2836
rect 4695 2787 5230 2821
rect 4695 2774 4704 2787
rect 5230 2772 5282 2778
rect 2380 2430 4490 2476
rect 1201 2304 1253 2310
rect 2380 2301 2426 2430
rect 3553 2304 3605 2310
rect 1253 2255 3553 2301
rect 1201 2246 1253 2252
rect 3553 2246 3605 2252
rect 1919 2122 1971 2128
rect 2835 2122 2887 2128
rect 1971 2073 2835 2119
rect 1919 2064 1971 2070
rect 613 1972 665 1978
rect 613 1914 665 1920
rect 622 1592 656 1914
rect 737 1867 743 1919
rect 795 1867 801 1919
rect 746 1592 792 1867
rect 613 1586 665 1592
rect 613 1528 665 1534
rect 743 1586 795 1592
rect 2380 1567 2426 2073
rect 2835 2064 2887 2070
rect 4005 1859 4011 1911
rect 4063 1859 4069 1911
rect 4014 1594 4060 1859
rect 4011 1588 4063 1594
rect 743 1528 795 1534
rect 2377 1561 2429 1567
rect 207 1424 572 1458
rect 746 1448 792 1528
rect 4011 1530 4063 1536
rect 2377 1503 2429 1509
rect 4014 1448 4060 1530
rect 155 1409 207 1415
rect 746 1402 4060 1448
rect 1032 450 1084 456
rect 1629 450 1681 456
rect 1084 401 1629 447
rect 1032 392 1084 398
rect 1919 450 1971 456
rect 1681 401 1919 447
rect 1629 392 1681 398
rect 2835 450 2887 456
rect 1971 401 2835 447
rect 1919 392 1971 398
rect 3127 450 3179 456
rect 2887 401 3127 447
rect 2835 392 2887 398
rect 3721 450 3773 456
rect 3179 401 3721 447
rect 3127 392 3179 398
rect 3721 392 3773 398
<< via2 >>
rect 4060 2774 4120 2834
rect 4635 2774 4695 2834
<< metal3 >>
rect 4055 2834 4125 2839
rect 4630 2834 4700 2839
rect 4055 2774 4060 2834
rect 4120 2774 4635 2834
rect 4695 2774 4700 2834
rect 4055 2769 4125 2774
rect 4630 2769 4700 2774
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_0
timestamp 1698929273
transform 1 0 998 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_1
timestamp 1698929273
transform 1 0 1586 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_2
timestamp 1698929273
transform 1 0 2174 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_3
timestamp 1698929273
transform 1 0 2632 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_4
timestamp 1698929273
transform 1 0 3220 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_5
timestamp 1698929273
transform 1 0 4396 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_6
timestamp 1698929273
transform 1 0 3220 0 1 1234
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_7
timestamp 1698929273
transform 1 0 1586 0 1 1234
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_8
timestamp 1698929273
transform 1 0 3808 0 1 1234
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_9
timestamp 1698929273
transform 1 0 410 0 1 1234
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_10
timestamp 1698929273
transform 1 0 998 0 1 1234
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_11
timestamp 1698929273
transform 1 0 -178 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_12
timestamp 1698929273
transform 1 0 3808 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CM22X2  sky130_fd_pr__nfet_g5v0d10v5_CM22X2_13
timestamp 1698929273
transform 1 0 410 0 1 2287
box -258 -457 258 457
use sky130_fd_pr__nfet_g5v0d10v5_CMVU23  sky130_fd_pr__nfet_g5v0d10v5_CMVU23_0
timestamp 1698929273
transform 1 0 2174 0 1 834
box -258 -857 258 857
use sky130_fd_pr__nfet_g5v0d10v5_CMVU23  sky130_fd_pr__nfet_g5v0d10v5_CMVU23_1
timestamp 1698929273
transform 1 0 -178 0 1 834
box -258 -857 258 857
use sky130_fd_pr__nfet_g5v0d10v5_CMVU23  sky130_fd_pr__nfet_g5v0d10v5_CMVU23_2
timestamp 1698929273
transform 1 0 4396 0 1 834
box -258 -857 258 857
use sky130_fd_pr__nfet_g5v0d10v5_CMVU23  sky130_fd_pr__nfet_g5v0d10v5_CMVU23_3
timestamp 1698929273
transform 1 0 2632 0 1 834
box -258 -857 258 857
use sky130_fd_pr__nfet_g5v0d10v5_JSTQTR  sky130_fd_pr__nfet_g5v0d10v5_JSTQTR_0
timestamp 1698929273
transform 1 0 5047 0 1 1354
box -108 -1377 108 1377
use sky130_fd_pr__nfet_g5v0d10v5_JSTQTR  sky130_fd_pr__nfet_g5v0d10v5_JSTQTR_1
timestamp 1698929273
transform 1 0 5623 0 1 1354
box -108 -1377 108 1377
use sky130_fd_pr__nfet_g5v0d10v5_JSTQTR  sky130_fd_pr__nfet_g5v0d10v5_JSTQTR_2
timestamp 1698929273
transform 1 0 5911 0 1 1354
box -108 -1377 108 1377
use sky130_fd_pr__nfet_g5v0d10v5_K5LT42  sky130_fd_pr__nfet_g5v0d10v5_K5LT42_0
timestamp 1698929273
transform 1 0 410 0 1 334
box -258 -357 258 357
use sky130_fd_pr__nfet_g5v0d10v5_KRRUZH  sky130_fd_pr__nfet_g5v0d10v5_KRRUZH_0
timestamp 1698929273
transform 1 0 5335 0 1 574
box -108 -597 108 597
use sky130_fd_pr__nfet_g5v0d10v5_NYRQZ6  sky130_fd_pr__nfet_g5v0d10v5_NYRQZ6_0
timestamp 1698929273
transform 1 0 5335 0 1 2487
box -108 -257 108 257
use sky130_fd_pr__nfet_g5v0d10v5_TNTUPH  sky130_fd_pr__nfet_g5v0d10v5_TNTUPH_1
timestamp 1698929273
transform 1 0 5335 0 1 1715
box -108 -457 108 457
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_0
timestamp 1698929273
transform 1 0 -178 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_2
timestamp 1698929273
transform 1 0 4396 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_3
timestamp 1698929273
transform 1 0 410 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_6
timestamp 1698929273
transform 1 0 998 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_7
timestamp 1698929273
transform 1 0 1586 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_8
timestamp 1698929273
transform 1 0 2174 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_9
timestamp 1698929273
transform 1 0 2632 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_10
timestamp 1698929273
transform 1 0 3220 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_EHRSHC  sky130_fd_pr__pfet_g5v0d10v5_EHRSHC_11
timestamp 1698929273
transform 1 0 3808 0 1 4186
box -324 -466 324 466
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_0
timestamp 1698929273
transform 1 0 -178 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_2
timestamp 1698929273
transform 1 0 4396 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_3
timestamp 1698929273
transform 1 0 410 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_6
timestamp 1698929273
transform 1 0 998 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_7
timestamp 1698929273
transform 1 0 1586 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_8
timestamp 1698929273
transform 1 0 3808 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_9
timestamp 1698929273
transform 1 0 3220 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_10
timestamp 1698929273
transform 1 0 2632 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_MBRSZA  sky130_fd_pr__pfet_g5v0d10v5_MBRSZA_11
timestamp 1698929273
transform 1 0 2174 0 1 3234
box -324 -364 324 402
use sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5  sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_0
timestamp 1698929273
transform 1 0 5623 0 1 3750
box -174 -864 174 902
use sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5  sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_1
timestamp 1698929273
transform 1 0 5911 0 1 3750
box -174 -864 174 902
use sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5  sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_2
timestamp 1698929273
transform 1 0 5335 0 1 3750
box -174 -864 174 902
use sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5  sky130_fd_pr__pfet_g5v0d10v5_UK4LZ5_3
timestamp 1698929273
transform 1 0 5047 0 1 3750
box -174 -864 174 902
use sky130_fd_pr__res_generic_nd__hv_USEA7F  sky130_fd_pr__res_generic_nd__hv_USEA7F_0
timestamp 1698929273
transform 1 0 3223 0 1 394
box -118 -346 118 348
use sky130_fd_pr__res_generic_nd__hv_USEA7F  sky130_fd_pr__res_generic_nd__hv_USEA7F_1
timestamp 1698929273
transform 1 0 1583 0 1 394
box -118 -346 118 348
use sky130_fd_pr__res_generic_nd__hv_USEA7F  sky130_fd_pr__res_generic_nd__hv_USEA7F_2
timestamp 1698929273
transform 1 0 3818 0 1 394
box -118 -346 118 348
use sky130_fd_pr__res_generic_nd__hv_USEA7F  sky130_fd_pr__res_generic_nd__hv_USEA7F_3
timestamp 1698929273
transform 1 0 988 0 1 394
box -118 -346 118 348
<< labels >>
flabel metal1 s 2996 -56 2996 -56 0 FreeSans 800 0 0 0 VSS
flabel metal1 s 2404 4676 2404 4676 0 FreeSans 800 0 0 0 VCC
flabel metal2 s 5193 2917 5193 2917 0 FreeSans 800 0 0 0 Vb2
flabel locali s 5539 2924 5539 2924 0 FreeSans 800 0 0 0 Vb1
flabel locali s 5257 2725 5257 2725 0 FreeSans 800 0 0 0 Vb3
flabel locali s 5416 2138 5416 2138 0 FreeSans 800 0 0 0 Vb5
<< end >>
