magic
tech sky130A
timestamp 1697281155
<< error_p >>
rect -87 -233 87 233
<< nwell >>
rect -72 -231 72 231
<< mvpmos >>
rect -25 -200 25 200
<< mvpdiff >>
rect -54 194 -25 200
rect -54 -194 -48 194
rect -31 -194 -25 194
rect -54 -200 -25 -194
rect 25 194 54 200
rect 25 -194 31 194
rect 48 -194 54 194
rect 25 -200 54 -194
<< mvpdiffc >>
rect -48 -194 -31 194
rect 31 -194 48 194
<< poly >>
rect -25 200 25 213
rect -25 -213 25 -200
<< locali >>
rect -48 194 -31 202
rect -48 -202 -31 -194
rect 31 194 48 202
rect 31 -202 48 -194
<< viali >>
rect -48 -194 -31 194
rect 31 -194 48 194
<< metal1 >>
rect -51 194 -28 200
rect -51 -194 -48 194
rect -31 -194 -28 194
rect -51 -200 -28 -194
rect 28 194 51 200
rect 28 -194 31 194
rect 48 -194 51 194
rect 28 -200 51 -194
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
