magic
tech sky130A
magscale 1 2
timestamp 1696698053
<< mvnmos >>
rect -300 -81 300 19
<< mvndiff >>
rect -358 7 -300 19
rect -358 -69 -346 7
rect -312 -69 -300 7
rect -358 -81 -300 -69
rect 300 7 358 19
rect 300 -69 312 7
rect 346 -69 358 7
rect 300 -81 358 -69
<< mvndiffc >>
rect -346 -69 -312 7
rect 312 -69 346 7
<< poly >>
rect -300 91 300 107
rect -300 57 -284 91
rect 284 57 300 91
rect -300 19 300 57
rect -300 -107 300 -81
<< polycont >>
rect -284 57 284 91
<< locali >>
rect -300 57 -284 91
rect 284 57 300 91
rect -346 7 -312 23
rect -346 -85 -312 -69
rect 312 7 346 23
rect 312 -85 346 -69
<< viali >>
rect -284 57 284 91
rect -346 -69 -312 7
rect 312 -69 346 7
<< metal1 >>
rect -296 91 296 97
rect -296 57 -284 91
rect 284 57 296 91
rect -296 51 296 57
rect -352 7 -306 19
rect -352 -69 -346 7
rect -312 -69 -306 7
rect -352 -81 -306 -69
rect 306 7 352 19
rect 306 -69 312 7
rect 346 -69 352 7
rect 306 -81 352 -69
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
