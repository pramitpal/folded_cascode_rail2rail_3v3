magic
tech sky130A
magscale 1 2
timestamp 1697281155
<< error_p >>
rect -144 430 144 464
rect -174 -502 174 430
<< nwell >>
rect -144 -498 144 464
<< mvpmos >>
rect -50 -436 50 364
<< mvpdiff >>
rect -108 352 -50 364
rect -108 -424 -96 352
rect -62 -424 -50 352
rect -108 -436 -50 -424
rect 50 352 108 364
rect 50 -424 62 352
rect 96 -424 108 352
rect 50 -436 108 -424
<< mvpdiffc >>
rect -96 -424 -62 352
rect 62 -424 96 352
<< poly >>
rect -50 445 50 461
rect -50 411 -34 445
rect 34 411 50 445
rect -50 364 50 411
rect -50 -462 50 -436
<< polycont >>
rect -34 411 34 445
<< locali >>
rect -50 411 -34 445
rect 34 411 50 445
rect -96 352 -62 368
rect -96 -440 -62 -424
rect 62 352 96 368
rect 62 -440 96 -424
<< viali >>
rect -34 411 34 445
rect -96 -424 -62 352
rect 62 -424 96 352
<< metal1 >>
rect -46 445 46 451
rect -46 411 -34 445
rect 34 411 46 445
rect -46 405 46 411
rect -102 352 -56 364
rect -102 -424 -96 352
rect -62 -424 -56 352
rect -102 -436 -56 -424
rect 56 352 102 364
rect 56 -424 62 352
rect 96 -424 102 352
rect 56 -436 102 -424
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
