magic
tech sky130A
magscale 1 2
timestamp 1698912251
<< mvnmos >>
rect -200 -381 200 319
<< mvndiff >>
rect -258 307 -200 319
rect -258 -369 -246 307
rect -212 -369 -200 307
rect -258 -381 -200 -369
rect 200 307 258 319
rect 200 -369 212 307
rect 246 -369 258 307
rect 200 -381 258 -369
<< mvndiffc >>
rect -246 -369 -212 307
rect 212 -369 246 307
<< poly >>
rect -200 391 200 407
rect -200 357 -184 391
rect 184 357 200 391
rect -200 319 200 357
rect -200 -407 200 -381
<< polycont >>
rect -184 357 184 391
<< locali >>
rect -200 357 -184 391
rect 184 357 200 391
rect -246 307 -212 323
rect -246 -385 -212 -369
rect 212 307 246 323
rect 212 -385 246 -369
<< viali >>
rect -184 357 184 391
rect -246 -369 -212 307
rect 212 -369 246 307
<< metal1 >>
rect -196 391 196 397
rect -196 357 -184 391
rect 184 357 196 391
rect -196 351 196 357
rect -252 307 -206 319
rect -252 -369 -246 307
rect -212 -369 -206 307
rect -252 -381 -206 -369
rect 206 307 252 319
rect 206 -369 212 307
rect 246 -369 252 307
rect 206 -381 252 -369
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.5 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
