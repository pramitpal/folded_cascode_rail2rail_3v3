magic
tech sky130A
magscale 1 2
timestamp 1697135688
<< nwell >>
rect -742 -343 1171 1100
<< mvpsubdiff >>
rect -670 -520 -622 -486
rect -670 -1866 -664 -520
rect -628 -1866 -622 -520
rect 1051 -520 1099 -486
rect -670 -1905 -622 -1866
rect 1051 -1866 1057 -520
rect 1093 -1866 1099 -520
rect 1051 -1905 1099 -1866
<< mvnsubdiff >>
rect -670 961 -622 1000
rect -670 -234 -664 961
rect -628 -234 -622 961
rect 1051 961 1099 1000
rect -670 -266 -622 -234
rect 1051 -234 1057 961
rect 1093 -234 1099 961
rect 1051 -266 1099 -234
<< mvpsubdiffcont >>
rect -664 -1866 -628 -520
rect 1057 -1866 1093 -520
<< mvnsubdiffcont >>
rect -664 -234 -628 961
rect 1057 -234 1093 961
<< poly >>
rect -202 153 -102 200
rect -202 119 -186 153
rect -118 119 -102 153
rect -202 103 -102 119
rect 86 153 186 200
rect 86 119 102 153
rect 170 119 186 153
rect 86 103 186 119
rect 244 153 344 200
rect 244 119 260 153
rect 328 119 344 153
rect 244 103 344 119
rect 532 153 632 200
rect 532 119 548 153
rect 616 119 632 153
rect 532 103 632 119
rect -202 15 -102 31
rect -202 -19 -186 15
rect -118 -19 -102 15
rect -202 -66 -102 -19
rect 86 15 186 31
rect 86 -19 102 15
rect 170 -19 186 15
rect 86 -66 186 -19
rect 244 15 344 31
rect 244 -19 260 15
rect 328 -19 344 15
rect 244 -66 344 -19
rect 532 15 632 31
rect 532 -19 548 15
rect 616 -19 632 15
rect 532 -66 632 -19
rect -202 -405 -102 -389
rect -202 -439 -186 -405
rect -118 -439 -102 -405
rect -202 -486 -102 -439
rect 86 -405 186 -389
rect 86 -439 102 -405
rect 170 -439 186 -405
rect 86 -486 186 -439
rect 244 -405 344 -389
rect 244 -439 260 -405
rect 328 -439 344 -405
rect 244 -486 344 -439
rect 532 -405 632 -389
rect 532 -439 548 -405
rect 616 -439 632 -405
rect 532 -486 632 -439
rect -202 -1024 -102 -1008
rect -202 -1058 -186 -1024
rect -118 -1058 -102 -1024
rect -202 -1105 -102 -1058
rect 86 -1024 186 -1008
rect 86 -1058 102 -1024
rect 170 -1058 186 -1024
rect 86 -1105 186 -1058
rect 244 -1024 344 -1008
rect 244 -1058 260 -1024
rect 328 -1058 344 -1024
rect 244 -1105 344 -1058
rect 532 -1024 632 -1008
rect 532 -1058 548 -1024
rect 616 -1058 632 -1024
rect 532 -1105 632 -1058
<< polycont >>
rect -186 119 -118 153
rect 102 119 170 153
rect 260 119 328 153
rect 548 119 616 153
rect -186 -19 -118 15
rect 102 -19 170 15
rect 260 -19 328 15
rect 548 -19 616 15
rect -186 -439 -118 -405
rect 102 -439 170 -405
rect 260 -439 328 -405
rect 548 -439 616 -405
rect -186 -1058 -118 -1024
rect 102 -1058 170 -1024
rect 260 -1058 328 -1024
rect 548 -1058 616 -1024
<< locali >>
rect -536 1047 966 1081
rect -670 988 -622 1000
rect -536 988 -502 1047
rect -670 961 -502 988
rect -670 -234 -664 961
rect -628 918 -502 961
rect -378 960 -344 1047
rect -247 986 -213 1047
rect 198 952 232 1047
rect 644 942 678 1047
rect 774 960 808 1047
rect 932 988 966 1047
rect 1051 988 1099 1000
rect 932 961 1099 988
rect -628 212 -531 918
rect 932 212 1057 961
rect -628 -78 -622 212
rect -202 119 -186 153
rect -118 119 102 153
rect 170 119 260 153
rect 328 119 548 153
rect 616 119 632 153
rect -16 50 446 84
rect -536 -19 -344 15
rect -202 -19 -186 15
rect -118 -19 102 15
rect 170 -19 260 15
rect 328 -19 548 15
rect 616 -19 632 15
rect 774 -19 966 15
rect -536 -78 -502 -19
rect -378 -78 -344 -19
rect -628 -122 -502 -78
rect 774 -103 808 -19
rect 932 -78 966 -19
rect 1051 -78 1057 212
rect -628 -234 -534 -122
rect -670 -254 -534 -234
rect 932 -234 1057 -78
rect 1093 -234 1099 961
rect 932 -254 1099 -234
rect -670 -266 -622 -254
rect 1051 -266 1099 -254
rect 93 -353 401 -319
rect -202 -439 -186 -405
rect -118 -439 102 -405
rect 170 -439 260 -405
rect 328 -439 548 -405
rect 616 -439 632 -405
rect -670 -520 -622 -486
rect 1051 -498 1099 -486
rect 931 -520 1099 -498
rect -670 -1866 -664 -520
rect -628 -857 -534 -520
rect -628 -874 -502 -857
rect -628 -1117 -622 -874
rect -536 -924 -502 -874
rect -378 -924 -344 -864
rect -536 -958 -344 -924
rect 773 -924 807 -862
rect 931 -874 1057 -520
rect 931 -924 965 -874
rect -10 -964 440 -930
rect 773 -958 965 -924
rect -202 -1058 -186 -1024
rect -118 -1058 102 -1024
rect 170 -1058 260 -1024
rect 328 -1058 548 -1024
rect 616 -1058 632 -1024
rect 1051 -1117 1057 -874
rect -628 -1866 -530 -1117
rect -670 -1874 -530 -1866
rect -670 -1893 -502 -1874
rect -670 -1905 -622 -1893
rect -536 -1943 -502 -1893
rect -378 -1943 -344 -1882
rect -248 -1943 -214 -1864
rect 931 -1866 1057 -1117
rect 1093 -1866 1099 -520
rect 198 -1943 232 -1891
rect 644 -1943 678 -1871
rect 773 -1943 807 -1884
rect 931 -1893 1099 -1866
rect 931 -1943 965 -1893
rect 1051 -1905 1099 -1893
rect -536 -1977 965 -1943
<< viali >>
rect -50 50 -16 84
rect 446 50 480 84
rect 59 -353 93 -319
rect 401 -353 435 -319
rect -44 -964 -10 -930
rect 440 -964 474 -930
<< metal1 >>
rect -90 96 -56 237
rect -90 84 -10 96
rect -90 50 -50 84
rect -16 50 -10 84
rect -90 38 -10 50
rect 40 84 74 226
rect 357 84 391 245
rect 486 96 520 242
rect 40 50 391 84
rect -248 -319 -214 -193
rect -90 -270 -56 38
rect 40 -254 74 50
rect 47 -319 105 -313
rect -248 -353 59 -319
rect 93 -353 105 -319
rect -248 -514 -214 -353
rect 47 -359 105 -353
rect 198 -533 232 -114
rect 357 -124 391 50
rect 440 84 520 96
rect 440 50 446 84
rect 480 50 520 84
rect 440 38 520 50
rect 486 -104 520 38
rect 389 -319 447 -313
rect 644 -319 678 -237
rect 389 -353 401 -319
rect 435 -353 678 -319
rect 389 -359 447 -353
rect 644 -560 678 -353
rect -90 -924 -56 -832
rect -90 -930 2 -924
rect -90 -964 -44 -930
rect -10 -964 2 -930
rect -90 -970 2 -964
rect 40 -930 74 -824
rect 356 -930 390 -800
rect 486 -924 520 -862
rect 40 -964 390 -930
rect -90 -1909 -56 -970
rect 40 -1893 74 -964
rect 356 -1893 390 -964
rect 428 -930 520 -924
rect 428 -964 440 -930
rect 474 -964 520 -930
rect 428 -970 520 -964
rect 486 -1909 520 -970
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_0
timestamp 1696962984
transform 1 0 294 0 1 -686
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_1
timestamp 1696962984
transform 1 0 582 0 1 -686
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_2
timestamp 1696962984
transform 1 0 136 0 1 -686
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_4
timestamp 1696962984
transform 1 0 -152 0 1 -686
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NYY6SB  sky130_fd_pr__nfet_g5v0d10v5_NYY6SB_0
timestamp 1696961404
transform 1 0 -440 0 1 -717
box -108 -257 108 257
use sky130_fd_pr__nfet_g5v0d10v5_NYY6SB  sky130_fd_pr__nfet_g5v0d10v5_NYY6SB_1
timestamp 1696961404
transform 1 0 869 0 1 -717
box -108 -257 108 257
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_0
timestamp 1696959484
transform 1 0 -152 0 1 -1505
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_1
timestamp 1696959484
transform 1 0 294 0 1 -1505
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_2
timestamp 1696959484
transform 1 0 136 0 1 -1505
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_3
timestamp 1696959484
transform 1 0 582 0 1 -1505
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNWANH  sky130_fd_pr__nfet_g5v0d10v5_TNWANH_0
timestamp 1696961404
transform 1 0 -440 0 1 -1536
box -108 -457 108 457
use sky130_fd_pr__nfet_g5v0d10v5_TNWANH  sky130_fd_pr__nfet_g5v0d10v5_TNWANH_1
timestamp 1696961404
transform 1 0 869 0 1 -1536
box -108 -457 108 457
use sky130_fd_pr__pfet_g5v0d10v5_DEERZ7  sky130_fd_pr__pfet_g5v0d10v5_DEERZ7_0
timestamp 1696961038
transform 1 0 -440 0 1 636
box -174 -502 174 464
use sky130_fd_pr__pfet_g5v0d10v5_DEERZ7  sky130_fd_pr__pfet_g5v0d10v5_DEERZ7_1
timestamp 1696961038
transform 1 0 870 0 1 636
box -174 -502 174 464
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_0
timestamp 1696958486
transform 1 0 -152 0 1 600
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_1
timestamp 1696958486
transform 1 0 136 0 1 600
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_2
timestamp 1696958486
transform 1 0 294 0 1 600
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_3
timestamp 1696958486
transform 1 0 582 0 1 600
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_0
timestamp 1696958827
transform 1 0 136 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_1
timestamp 1696958827
transform 1 0 -152 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_2
timestamp 1696958827
transform 1 0 294 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_3
timestamp 1696958827
transform 1 0 582 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7  sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_0
timestamp 1696961150
transform 1 0 -440 0 1 -130
box -174 -202 174 164
use sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7  sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_1
timestamp 1696961150
transform 1 0 870 0 1 -130
box -174 -202 174 164
<< labels >>
flabel locali s 212 1066 212 1066 0 FreeSans 800 0 0 0 VCC
flabel locali s 214 -1955 214 -1955 0 FreeSans 800 0 0 0 VSS
flabel locali s 442 -1034 442 -1034 0 FreeSans 800 0 0 0 CMFB
flabel locali s 437 -425 437 -425 0 FreeSans 800 0 0 0 Vb3
flabel locali s 442 2 442 2 0 FreeSans 800 0 0 0 Vb2
flabel locali s 440 138 440 138 0 FreeSans 800 0 0 0 Vb1
flabel metal1 s 219 -381 219 -381 0 FreeSans 800 0 0 0 out
flabel metal1 s 663 -381 663 -381 0 FreeSans 800 0 0 0 out2
flabel metal1 s 57 96 57 96 0 FreeSans 800 0 0 0 N2
flabel metal1 s -75 35 -75 35 0 FreeSans 800 0 0 0 N1
flabel metal1 s 56 -987 56 -987 0 FreeSans 800 0 0 0 N4
flabel metal1 s -75 -1083 -75 -1083 0 FreeSans 800 0 0 0 N3
<< end >>
