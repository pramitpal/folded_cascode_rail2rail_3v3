magic
tech sky130A
magscale 1 2
timestamp 1697289488
<< error_p >>
rect -144 830 144 864
rect -174 -902 174 830
<< nwell >>
rect -144 -898 144 864
<< mvpmos >>
rect -50 -836 50 764
<< mvpdiff >>
rect -108 752 -50 764
rect -108 -824 -96 752
rect -62 -824 -50 752
rect -108 -836 -50 -824
rect 50 752 108 764
rect 50 -824 62 752
rect 96 -824 108 752
rect 50 -836 108 -824
<< mvpdiffc >>
rect -96 -824 -62 752
rect 62 -824 96 752
<< poly >>
rect -50 845 50 861
rect -50 811 -34 845
rect 34 811 50 845
rect -50 764 50 811
rect -50 -862 50 -836
<< polycont >>
rect -34 811 34 845
<< locali >>
rect -50 811 -34 845
rect 34 811 50 845
rect -96 752 -62 768
rect -96 -840 -62 -824
rect 62 752 96 768
rect 62 -840 96 -824
<< viali >>
rect -34 811 34 845
rect -96 -824 -62 752
rect 62 -824 96 752
<< metal1 >>
rect -46 845 46 851
rect -46 811 -34 845
rect 34 811 46 845
rect -46 805 46 811
rect -102 752 -56 764
rect -102 -824 -96 752
rect -62 -824 -56 752
rect -102 -836 -56 -824
rect 56 752 102 764
rect 56 -824 62 752
rect 96 -824 102 752
rect 56 -836 102 -824
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
