magic
tech sky130A
magscale 1 2
timestamp 1697289488
<< error_p >>
rect -108 -169 -50 231
rect 50 -169 108 231
<< mvnmos >>
rect -50 -169 50 231
<< mvndiff >>
rect -108 219 -50 231
rect -108 -157 -96 219
rect -62 -157 -50 219
rect -108 -169 -50 -157
rect 50 219 108 231
rect 50 -157 62 219
rect 96 -157 108 219
rect 50 -169 108 -157
<< mvndiffc >>
rect -96 -157 -62 219
rect 62 -157 96 219
<< poly >>
rect -50 231 50 257
rect -50 -207 50 -169
rect -50 -241 -34 -207
rect 34 -241 50 -207
rect -50 -257 50 -241
<< polycont >>
rect -34 -241 34 -207
<< locali >>
rect -96 219 -62 235
rect -96 -173 -62 -157
rect 62 219 96 235
rect 62 -173 96 -157
rect -50 -241 -34 -207
rect 34 -241 50 -207
<< viali >>
rect -96 -157 -62 219
rect 62 -157 96 219
rect -34 -241 34 -207
<< metal1 >>
rect -102 219 -56 231
rect -102 -157 -96 219
rect -62 -157 -56 219
rect -102 -169 -56 -157
rect 56 219 102 231
rect 56 -157 62 219
rect 96 -157 102 219
rect 56 -169 102 -157
rect -46 -207 46 -201
rect -46 -241 -34 -207
rect 34 -241 46 -207
rect -46 -247 46 -241
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
