magic
tech sky130A
timestamp 1698929273
<< error_p >>
rect -87 -58 87 58
<< nwell >>
rect -72 -56 72 56
<< mvpmos >>
rect -25 -25 25 25
<< mvpdiff >>
rect -54 19 -25 25
rect -54 -19 -48 19
rect -31 -19 -25 19
rect -54 -25 -25 -19
rect 25 19 54 25
rect 25 -19 31 19
rect 48 -19 54 19
rect 25 -25 54 -19
<< mvpdiffc >>
rect -48 -19 -31 19
rect 31 -19 48 19
<< poly >>
rect -25 25 25 38
rect -25 -38 25 -25
<< locali >>
rect -48 19 -31 27
rect -48 -27 -31 -19
rect 31 19 48 27
rect 31 -27 48 -19
<< viali >>
rect -48 -19 -31 19
rect 31 -19 48 19
<< metal1 >>
rect -51 19 -28 25
rect -51 -19 -48 19
rect -31 -19 -28 19
rect -51 -25 -28 -19
rect 28 19 51 25
rect 28 -19 31 19
rect 48 -19 51 19
rect 28 -25 51 -19
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
