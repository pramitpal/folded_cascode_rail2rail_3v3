magic
tech sky130A
timestamp 1697284980
<< error_p >>
rect -87 331 87 333
rect -87 -331 -72 331
rect -54 298 54 300
rect -54 -298 -39 298
rect 39 -298 54 298
rect -54 -300 54 -298
rect 72 -331 87 331
rect -87 -333 87 -331
<< nwell >>
rect -72 -331 72 331
<< mvpmos >>
rect -25 -300 25 300
<< mvpdiff >>
rect -54 294 -25 300
rect -54 -294 -48 294
rect -31 -294 -25 294
rect -54 -300 -25 -294
rect 25 294 54 300
rect 25 -294 31 294
rect 48 -294 54 294
rect 25 -300 54 -294
<< mvpdiffc >>
rect -48 -294 -31 294
rect 31 -294 48 294
<< poly >>
rect -25 300 25 313
rect -25 -313 25 -300
<< locali >>
rect -48 294 -31 302
rect -48 -302 -31 -294
rect 31 294 48 302
rect 31 -302 48 -294
<< viali >>
rect -48 -294 -31 294
rect 31 -294 48 294
<< metal1 >>
rect -51 294 -28 300
rect -51 -294 -48 294
rect -31 -294 -28 294
rect -51 -300 -28 -294
rect 28 294 51 300
rect 28 -294 31 294
rect 48 -294 51 294
rect 28 -300 51 -294
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
