magic
tech sky130A
magscale 1 2
timestamp 1698929273
<< error_p >>
rect -108 -571 -50 509
rect 50 -571 108 509
<< mvnmos >>
rect -50 -571 50 509
<< mvndiff >>
rect -108 497 -50 509
rect -108 -559 -96 497
rect -62 -559 -50 497
rect -108 -571 -50 -559
rect 50 497 108 509
rect 50 -559 62 497
rect 96 -559 108 497
rect 50 -571 108 -559
<< mvndiffc >>
rect -96 -559 -62 497
rect 62 -559 96 497
<< poly >>
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 509 50 547
rect -50 -597 50 -571
<< polycont >>
rect -34 547 34 581
<< locali >>
rect -50 547 -34 581
rect 34 547 50 581
rect -96 497 -62 513
rect -96 -575 -62 -559
rect 62 497 96 513
rect 62 -575 96 -559
<< viali >>
rect -34 547 34 581
rect -96 -559 -62 497
rect 62 -559 96 497
<< metal1 >>
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect -102 497 -56 509
rect -102 -559 -96 497
rect -62 -559 -56 497
rect -102 -571 -56 -559
rect 56 497 102 509
rect 56 -559 62 497
rect 96 -559 102 497
rect 56 -571 102 -559
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.4 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
