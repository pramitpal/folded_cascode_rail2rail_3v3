** sch_path:
*+ /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/backup_schematic/current_source.sch
.subckt current_source VCC VSS Vb1 Vb2 Vb3 Vb5
*.PININFO VCC:B VSS:B Vb1:O Vb2:O Vb3:O Vb5:O
XM23 Vb1 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM24 Vb2 Vb2 Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM25 Vb5 Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM26 Vb3 Vb3 Vb5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM58 net6 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM59 net1 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM60 net7 net4 net5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=4
XM61 net4 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM64 net2 net3 net6 VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 m=2
XM65 net3 net3 net1 VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 m=2
XM66 net3 net2 net7 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM67 net2 net2 net4 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM68 net8 net2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=2 nf=1 m=1
XM69 net8 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=1
XM70 net1 net8 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=2 nf=1 m=1
XM71 net9 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM72 Vb3 net3 net9 VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 m=2
XM73 net10 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM74 Vb2 net2 net10 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM11 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM12 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM13 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM14 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM15 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM16 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XR1 VSS net5 VSS sky130_fd_pr__res_generic_nd__hv W=0.42 L=6.927 mult=4 m=4
XM17 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM6 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM7 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM8 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM9 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM10 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM2 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM3 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM4 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
.ends
.end
