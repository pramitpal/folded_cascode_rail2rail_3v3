magic
tech sky130A
magscale 1 2
timestamp 1697281155
<< nwell >>
rect -742 -343 1171 1176
<< mvpsubdiff >>
rect -670 -590 -622 -556
rect -670 -2006 -664 -590
rect -628 -2006 -622 -590
rect 1051 -590 1099 -556
rect -670 -2045 -622 -2006
rect 1051 -2006 1057 -590
rect 1093 -2006 1099 -590
rect 1051 -2045 1099 -2006
<< mvnsubdiff >>
rect -670 1037 -622 1076
rect -670 -234 -664 1037
rect -628 -234 -622 1037
rect 1051 1037 1099 1076
rect -670 -266 -622 -234
rect 1051 -234 1057 1037
rect 1093 -234 1099 1037
rect 1051 -266 1099 -234
<< mvpsubdiffcont >>
rect -664 -2006 -628 -590
rect 1057 -2006 1093 -590
<< mvnsubdiffcont >>
rect -664 -234 -628 1037
rect 1057 -234 1093 1037
<< poly >>
rect -202 229 -102 276
rect -202 195 -186 229
rect -118 195 -102 229
rect -202 179 -102 195
rect 86 229 186 276
rect 86 195 102 229
rect 170 195 186 229
rect 86 179 186 195
rect 244 229 344 276
rect 244 195 260 229
rect 328 195 344 229
rect 244 179 344 195
rect 532 229 632 276
rect 532 195 548 229
rect 616 195 632 229
rect 532 179 632 195
rect -202 15 -102 31
rect -202 -19 -186 15
rect -118 -19 -102 15
rect -202 -66 -102 -19
rect 86 15 186 31
rect 86 -19 102 15
rect 170 -19 186 15
rect 86 -66 186 -19
rect 244 15 344 31
rect 244 -19 260 15
rect 328 -19 344 15
rect 244 -66 344 -19
rect 532 15 632 31
rect 532 -19 548 15
rect 616 -19 632 15
rect 532 -66 632 -19
rect -202 -475 -102 -459
rect -202 -509 -186 -475
rect -118 -509 -102 -475
rect -202 -556 -102 -509
rect 86 -475 186 -459
rect 86 -509 102 -475
rect 170 -509 186 -475
rect 86 -556 186 -509
rect 244 -475 344 -459
rect 244 -509 260 -475
rect 328 -509 344 -475
rect 244 -556 344 -509
rect 532 -475 632 -459
rect 532 -509 548 -475
rect 616 -509 632 -475
rect 532 -556 632 -509
rect -202 -1164 -102 -1148
rect -202 -1198 -186 -1164
rect -118 -1198 -102 -1164
rect -202 -1245 -102 -1198
rect 86 -1164 186 -1148
rect 86 -1198 102 -1164
rect 170 -1198 186 -1164
rect 86 -1245 186 -1198
rect 244 -1164 344 -1148
rect 244 -1198 260 -1164
rect 328 -1198 344 -1164
rect 244 -1245 344 -1198
rect 532 -1164 632 -1148
rect 532 -1198 548 -1164
rect 616 -1198 632 -1164
rect 532 -1245 632 -1198
<< polycont >>
rect -186 195 -118 229
rect 102 195 170 229
rect 260 195 328 229
rect 548 195 616 229
rect -186 -19 -118 15
rect 102 -19 170 15
rect 260 -19 328 15
rect 548 -19 616 15
rect -186 -509 -118 -475
rect 102 -509 170 -475
rect 260 -509 328 -475
rect 548 -509 616 -475
rect -186 -1198 -118 -1164
rect 102 -1198 170 -1164
rect 260 -1198 328 -1164
rect 548 -1198 616 -1164
<< locali >>
rect -536 1123 966 1157
rect -670 1064 -622 1076
rect -536 1064 -502 1123
rect -670 1037 -502 1064
rect -670 -234 -664 1037
rect -628 994 -502 1037
rect -378 1036 -344 1123
rect -247 1062 -213 1123
rect 198 1028 232 1123
rect 644 1018 678 1123
rect 774 1036 808 1123
rect 932 1064 966 1123
rect 1051 1064 1099 1076
rect 932 1037 1099 1064
rect -628 288 -531 994
rect 932 288 1057 1037
rect -628 -78 -622 288
rect -402 195 -186 229
rect -118 195 102 229
rect 170 195 260 229
rect 328 195 548 229
rect 616 195 632 229
rect -16 126 446 160
rect 198 86 232 126
rect -551 52 232 86
rect -536 -19 -344 15
rect -257 -19 -186 15
rect -118 -19 102 15
rect 170 -19 260 15
rect 328 -19 548 15
rect 616 -19 632 15
rect 774 -19 966 15
rect -536 -78 -502 -19
rect -378 -78 -344 -19
rect -628 -122 -502 -78
rect 774 -103 808 -19
rect 932 -78 966 -19
rect 1051 -78 1057 288
rect -628 -234 -534 -122
rect -670 -254 -534 -234
rect 932 -234 1057 -78
rect 1093 -234 1099 1037
rect 932 -254 1099 -234
rect -670 -266 -622 -254
rect 1051 -266 1099 -254
rect 93 -353 401 -319
rect 199 -396 233 -353
rect 199 -430 963 -396
rect -202 -509 -186 -475
rect -118 -509 102 -475
rect 170 -509 260 -475
rect 328 -509 548 -475
rect 616 -509 632 -475
rect -670 -590 -622 -556
rect 1051 -568 1099 -556
rect 931 -590 1099 -568
rect -670 -2006 -664 -590
rect -628 -927 -534 -590
rect -628 -944 -502 -927
rect -628 -1257 -622 -944
rect -536 -994 -502 -944
rect -378 -994 -344 -934
rect -536 -1028 -344 -994
rect 773 -994 807 -932
rect 931 -944 1057 -590
rect 931 -994 965 -944
rect -10 -1034 440 -1000
rect 773 -1028 965 -994
rect 198 -1073 232 -1034
rect -224 -1107 232 -1073
rect -202 -1198 -186 -1164
rect -118 -1198 102 -1164
rect 170 -1198 260 -1164
rect 328 -1198 548 -1164
rect 616 -1198 843 -1164
rect 1051 -1257 1057 -944
rect -628 -2006 -530 -1257
rect -670 -2014 -530 -2006
rect -670 -2033 -502 -2014
rect -670 -2045 -622 -2033
rect -536 -2083 -502 -2033
rect -378 -2083 -344 -2022
rect -248 -2083 -214 -2004
rect 931 -2006 1057 -1257
rect 1093 -2006 1099 -590
rect 198 -2083 232 -2031
rect 644 -2083 678 -2011
rect 773 -2083 807 -2024
rect 931 -2033 1099 -2006
rect 931 -2083 965 -2033
rect 1051 -2045 1099 -2033
rect -536 -2117 965 -2083
<< viali >>
rect -436 195 -402 229
rect -50 126 -16 160
rect 446 126 480 160
rect -585 52 -551 86
rect -291 -19 -257 15
rect 59 -353 93 -319
rect 401 -353 435 -319
rect -44 -1034 -10 -1000
rect 440 -1034 474 -1000
rect -258 -1107 -224 -1073
rect 843 -1198 877 -1164
<< metal1 >>
rect -442 229 -396 241
rect -742 195 -436 229
rect -402 195 -396 229
rect -442 183 -396 195
rect -90 172 -56 313
rect -351 120 -345 172
rect -293 163 -287 172
rect -293 120 -257 163
rect -591 86 -545 98
rect -742 52 -585 86
rect -551 52 -545 86
rect -591 40 -545 52
rect -291 27 -257 120
rect -90 160 -10 172
rect -90 126 -50 160
rect -16 126 -10 160
rect -90 114 -10 126
rect 40 160 74 302
rect 357 160 391 321
rect 486 172 520 318
rect 40 126 391 160
rect -297 15 -251 27
rect -297 -19 -291 15
rect -257 -19 -251 15
rect -297 -31 -251 -19
rect -248 -319 -214 -193
rect -90 -270 -56 114
rect 40 -254 74 126
rect 103 43 109 95
rect 161 86 167 95
rect 198 86 232 126
rect 161 52 232 86
rect 161 43 167 52
rect 47 -319 105 -313
rect -248 -353 59 -319
rect 93 -353 105 -319
rect -248 -584 -214 -353
rect 47 -359 105 -353
rect 198 -396 232 -114
rect 357 -124 391 126
rect 440 160 520 172
rect 440 126 446 160
rect 480 126 520 160
rect 440 114 520 126
rect 486 -104 520 114
rect 389 -319 447 -313
rect 644 -319 678 -237
rect 389 -353 401 -319
rect 435 -353 678 -319
rect 389 -359 447 -353
rect 533 -396 539 -387
rect 198 -430 539 -396
rect 198 -603 232 -430
rect 533 -439 539 -430
rect 591 -439 597 -387
rect 644 -630 678 -353
rect -90 -994 -56 -902
rect -90 -1000 2 -994
rect -90 -1034 -44 -1000
rect -10 -1034 2 -1000
rect -90 -1040 2 -1034
rect 40 -1000 74 -894
rect 356 -1000 390 -870
rect 486 -994 520 -932
rect 40 -1034 390 -1000
rect -264 -1073 -218 -1061
rect -327 -1107 -258 -1073
rect -224 -1107 -218 -1073
rect -264 -1119 -218 -1107
rect -90 -2049 -56 -1040
rect 40 -2033 74 -1034
rect 104 -1116 110 -1064
rect 162 -1073 168 -1064
rect 198 -1073 232 -1034
rect 162 -1107 232 -1073
rect 162 -1116 168 -1107
rect 356 -2033 390 -1034
rect 428 -1000 520 -994
rect 428 -1034 440 -1000
rect 474 -1034 520 -1000
rect 428 -1040 520 -1034
rect 486 -2049 520 -1040
rect 837 -1164 883 -1152
rect 837 -1198 843 -1164
rect 877 -1198 1199 -1164
rect 837 -1210 883 -1198
<< via1 >>
rect -345 120 -293 172
rect 109 43 161 95
rect 539 -439 591 -387
rect 110 -1116 162 -1064
<< metal2 >>
rect -345 172 -293 178
rect -742 129 -345 163
rect -345 114 -293 120
rect 109 95 161 101
rect -471 52 109 86
rect 109 37 161 43
rect 539 -387 591 -381
rect 591 -430 858 -396
rect 539 -445 591 -439
rect 110 -1064 162 -1058
rect -150 -1107 110 -1073
rect 110 -1122 162 -1116
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_0
timestamp 1697281155
transform 1 0 294 0 1 -756
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_1
timestamp 1697281155
transform 1 0 582 0 1 -756
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_2
timestamp 1697281155
transform 1 0 136 0 1 -756
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6#0  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_4
timestamp 1697281155
transform 1 0 -152 0 1 -756
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NYY6SB  sky130_fd_pr__nfet_g5v0d10v5_NYY6SB_0
timestamp 1697281155
transform 1 0 -440 0 1 -787
box -108 -257 108 257
use sky130_fd_pr__nfet_g5v0d10v5_NYY6SB  sky130_fd_pr__nfet_g5v0d10v5_NYY6SB_1
timestamp 1697281155
transform 1 0 869 0 1 -787
box -108 -257 108 257
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_0
timestamp 1697281155
transform 1 0 -152 0 1 -1645
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_1
timestamp 1697281155
transform 1 0 294 0 1 -1645
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_2
timestamp 1697281155
transform 1 0 136 0 1 -1645
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_3
timestamp 1697281155
transform 1 0 582 0 1 -1645
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_TNWANH  sky130_fd_pr__nfet_g5v0d10v5_TNWANH_0
timestamp 1697281155
transform 1 0 -440 0 1 -1676
box -108 -457 108 457
use sky130_fd_pr__nfet_g5v0d10v5_TNWANH  sky130_fd_pr__nfet_g5v0d10v5_TNWANH_1
timestamp 1697281155
transform 1 0 869 0 1 -1676
box -108 -457 108 457
use sky130_fd_pr__pfet_g5v0d10v5_DEERZ7  sky130_fd_pr__pfet_g5v0d10v5_DEERZ7_0
timestamp 1697281155
transform 1 0 -440 0 1 712
box -174 -502 174 464
use sky130_fd_pr__pfet_g5v0d10v5_DEERZ7  sky130_fd_pr__pfet_g5v0d10v5_DEERZ7_1
timestamp 1697281155
transform 1 0 870 0 1 712
box -174 -502 174 464
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_0
timestamp 1697281155
transform 1 0 -152 0 1 676
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_1
timestamp 1697281155
transform 1 0 136 0 1 676
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_2
timestamp 1697281155
transform 1 0 294 0 1 676
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_JEERZ7#0  sky130_fd_pr__pfet_g5v0d10v5_JEERZ7_3
timestamp 1697281155
transform 1 0 582 0 1 676
box -174 -466 174 466
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_0
timestamp 1697281155
transform 1 0 136 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_1
timestamp 1697281155
transform 1 0 -152 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_2
timestamp 1697281155
transform 1 0 294 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_3
timestamp 1697281155
transform 1 0 582 0 1 -166
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7  sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_0
timestamp 1697281155
transform 1 0 -440 0 1 -130
box -174 -202 174 164
use sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7  sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_1
timestamp 1697281155
transform 1 0 870 0 1 -130
box -174 -202 174 164
<< labels >>
flabel locali s 442 2 442 2 0 FreeSans 800 0 0 0 Vb2
flabel locali s 212 1142 212 1142 0 FreeSans 800 0 0 0 VCC
flabel locali s 440 214 440 214 0 FreeSans 800 0 0 0 Vb1
flabel metal1 s 57 172 57 172 0 FreeSans 800 0 0 0 N2
flabel metal1 s -75 111 -75 111 0 FreeSans 800 0 0 0 N1
flabel locali s 437 -495 437 -495 0 FreeSans 800 0 0 0 Vb3
flabel metal1 s 219 -451 219 -451 0 FreeSans 800 0 0 0 out
flabel metal1 s 663 -451 663 -451 0 FreeSans 800 0 0 0 out2
flabel metal1 s -75 -1223 -75 -1223 0 FreeSans 800 0 0 0 N3
flabel locali s 442 -1174 442 -1174 0 FreeSans 800 0 0 0 CMFB
flabel locali s 214 -2095 214 -2095 0 FreeSans 800 0 0 0 VSS
flabel metal1 s 56 -1061 56 -1061 0 FreeSans 800 0 0 0 N4
<< end >>
