** sch_path:
*+ /foss/designs/Comparator/old/schematic/folded_cascode/latest_working_comparator/backup_schematic/folded_cascode.sch
.subckt total VCC VSS INN INP VOUT
*.PININFO VCC:B VSS:B INN:I INP:I VOUT:O
XM23 Vb1 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM24 Vb2 Vb2 Vb1 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM25 Vb5 Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM26 Vb3 Vb3 Vb5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM58 net6 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM59 net1 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM60 net7 net4 net5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=4
XM61 net4 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM64 net2 net3 net6 VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 m=2
XM65 net3 net3 net1 VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 m=2
XM66 net3 net2 net7 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM67 net2 net2 net4 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM68 net8 net2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=2 nf=1 m=1
XM69 net8 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=1
XM70 net1 net8 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=2 nf=1 m=1
XM71 net9 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM72 Vb3 net3 net9 VCC sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 m=2
XM73 net17 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM74 Vb2 net2 net17 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4 nf=1 m=2
XM62 N2 INN net10 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM63 N1 INP net10 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM75 N3 INP net11 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM76 net11 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=4
XM77 net10 Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=4
XM78 N4 INN net11 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=2
XM79 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM80 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM81 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM82 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM83 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
XM84 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
XM85 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
XM86 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.5 nf=1 m=1
XM87 N4 CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=4
XM88 out Vb3 N4 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=4
XM89 out2 Vb3 N3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=4
XM90 N3 CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=4
XM91 out2 Vb2 N1 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=4
XM92 out Vb2 N2 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=4
XM93 N1 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=4
XM94 N2 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=4
XM95 VCC VCC VREF VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM96 VREF VREF VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM97 net12 net12 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.5 nf=1 m=2
XM98 v net12 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.5 nf=1 m=2
XM99 v out2 net13 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM100 net12 out net13 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM101 net13 Vb5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=4
XM102 VV v VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=6 nf=1 m=1
XM103 VV v VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM104 VOUT VV VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM105 VOUT VV VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM106 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=2 nf=1 m=1
XM107 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=0.5 nf=1 m=1
XM108 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=0.5 nf=1 m=1
XM109 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=2 nf=1 m=1
XM110 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM111 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM112 CMFB VREF net15 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=2
XM113 CMFB VREF net16 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=2
XM114 net14 out net15 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=2
XM115 net14 out2 net16 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=2
XM116 net15 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=2
XM117 net16 Vb1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=2
XM118 CMFB CMFB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.5 nf=1 m=2
XM119 net14 net14 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.5 nf=1 m=2
XM120 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.5 nf=1 m=1
XM121 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.5 nf=1 m=1
XM122 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM123 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM124 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM125 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM126 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM127 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM128 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM129 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM130 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM131 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM132 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM133 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XC1 CMFB VSS sky130_fd_pr__cap_mim_m3_1 W=7.1 L=6 m=1
XM11 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM12 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM13 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM14 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM15 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM16 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XR1 VSS net5 VSS sky130_fd_pr__res_generic_nd__hv W=0.42 L=6.927 mult=4 m=4
XM17 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM6 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM7 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM8 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM9 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM10 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM1 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM2 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM3 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
XM4 VCC VCC VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=1 m=1
.ends
.end
