magic
tech sky130A
magscale 1 2
timestamp 1697133871
<< mvnmos >>
rect -50 -19 50 81
<< mvndiff >>
rect -108 69 -50 81
rect -108 -7 -96 69
rect -62 -7 -50 69
rect -108 -19 -50 -7
rect 50 69 108 81
rect 50 -7 62 69
rect 96 -7 108 69
rect 50 -19 108 -7
<< mvndiffc >>
rect -96 -7 -62 69
rect 62 -7 96 69
<< poly >>
rect -50 81 50 107
rect -50 -57 50 -19
rect -50 -91 -34 -57
rect 34 -91 50 -57
rect -50 -107 50 -91
<< polycont >>
rect -34 -91 34 -57
<< locali >>
rect -96 69 -62 85
rect -96 -23 -62 -7
rect 62 69 96 85
rect 62 -23 96 -7
rect -50 -91 -34 -57
rect 34 -91 50 -57
<< viali >>
rect -96 -7 -62 69
rect 62 -7 96 69
rect -34 -91 34 -57
<< metal1 >>
rect -102 69 -56 81
rect -102 -7 -96 69
rect -62 -7 -56 69
rect -102 -19 -56 -7
rect 56 69 102 81
rect 56 -7 62 69
rect 96 -7 102 69
rect 56 -19 102 -7
rect -46 -57 46 -51
rect -46 -91 -34 -57
rect 34 -91 46 -57
rect -46 -97 46 -91
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
