magic
tech sky130A
timestamp 1697286120
<< error_p >>
rect -87 531 87 533
rect -87 -531 -72 531
rect -54 498 54 500
rect -54 -498 -39 498
rect 39 -498 54 498
rect -54 -500 54 -498
rect 72 -531 87 531
rect -87 -533 87 -531
<< nwell >>
rect -72 -531 72 531
<< mvpmos >>
rect -25 -500 25 500
<< mvpdiff >>
rect -54 494 -25 500
rect -54 -494 -48 494
rect -31 -494 -25 494
rect -54 -500 -25 -494
rect 25 494 54 500
rect 25 -494 31 494
rect 48 -494 54 494
rect 25 -500 54 -494
<< mvpdiffc >>
rect -48 -494 -31 494
rect 31 -494 48 494
<< poly >>
rect -25 500 25 513
rect -25 -513 25 -500
<< locali >>
rect -48 494 -31 502
rect -48 -502 -31 -494
rect 31 494 48 502
rect 31 -502 48 -494
<< viali >>
rect -48 -494 -31 494
rect 31 -494 48 494
<< metal1 >>
rect -51 494 -28 500
rect -51 -494 -48 494
rect -31 -494 -28 494
rect -51 -500 -28 -494
rect 28 494 51 500
rect 28 -494 31 494
rect 48 -494 51 494
rect 28 -500 51 -494
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
