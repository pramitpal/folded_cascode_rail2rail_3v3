magic
tech sky130A
magscale 1 2
timestamp 1698929273
<< error_p >>
rect -108 -769 -50 831
rect 50 -769 108 831
<< mvnmos >>
rect -50 -769 50 831
<< mvndiff >>
rect -108 819 -50 831
rect -108 -757 -96 819
rect -62 -757 -50 819
rect -108 -769 -50 -757
rect 50 819 108 831
rect 50 -757 62 819
rect 96 -757 108 819
rect 50 -769 108 -757
<< mvndiffc >>
rect -96 -757 -62 819
rect 62 -757 96 819
<< poly >>
rect -50 831 50 857
rect -50 -807 50 -769
rect -50 -841 -34 -807
rect 34 -841 50 -807
rect -50 -857 50 -841
<< polycont >>
rect -34 -841 34 -807
<< locali >>
rect -96 819 -62 835
rect -96 -773 -62 -757
rect 62 819 96 835
rect 62 -773 96 -757
rect -50 -841 -34 -807
rect 34 -841 50 -807
<< viali >>
rect -96 -757 -62 819
rect 62 -757 96 819
rect -34 -841 34 -807
<< metal1 >>
rect -102 819 -56 831
rect -102 -757 -96 819
rect -62 -757 -56 819
rect -102 -769 -56 -757
rect 56 819 102 831
rect 56 -757 62 819
rect 96 -757 102 819
rect 56 -769 102 -757
rect -46 -807 46 -801
rect -46 -841 -34 -807
rect 34 -841 46 -807
rect -46 -847 46 -841
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
