magic
tech sky130A
magscale 1 2
timestamp 1698695308
<< xpolycontact >>
rect -616 250 -546 682
rect -616 -682 -546 -250
rect -450 250 -380 682
rect -450 -682 -380 -250
rect -284 250 -214 682
rect -284 -682 -214 -250
rect -118 250 -48 682
rect -118 -682 -48 -250
rect 48 250 118 682
rect 48 -682 118 -250
rect 214 250 284 682
rect 214 -682 284 -250
rect 380 250 450 682
rect 380 -682 450 -250
rect 546 250 616 682
rect 546 -682 616 -250
<< ppolyres >>
rect -616 -250 -546 250
rect -450 -250 -380 250
rect -284 -250 -214 250
rect -118 -250 -48 250
rect 48 -250 118 250
rect 214 -250 284 250
rect 380 -250 450 250
rect 546 -250 616 250
<< viali >>
rect -600 267 -562 664
rect -434 267 -396 664
rect -268 267 -230 664
rect -102 267 -64 664
rect 64 267 102 664
rect 230 267 268 664
rect 396 267 434 664
rect 562 267 600 664
rect -600 -664 -562 -267
rect -434 -664 -396 -267
rect -268 -664 -230 -267
rect -102 -664 -64 -267
rect 64 -664 102 -267
rect 230 -664 268 -267
rect 396 -664 434 -267
rect 562 -664 600 -267
<< metal1 >>
rect -606 664 -556 676
rect -606 267 -600 664
rect -562 267 -556 664
rect -606 255 -556 267
rect -440 664 -390 676
rect -440 267 -434 664
rect -396 267 -390 664
rect -440 255 -390 267
rect -274 664 -224 676
rect -274 267 -268 664
rect -230 267 -224 664
rect -274 255 -224 267
rect -108 664 -58 676
rect -108 267 -102 664
rect -64 267 -58 664
rect -108 255 -58 267
rect 58 664 108 676
rect 58 267 64 664
rect 102 267 108 664
rect 58 255 108 267
rect 224 664 274 676
rect 224 267 230 664
rect 268 267 274 664
rect 224 255 274 267
rect 390 664 440 676
rect 390 267 396 664
rect 434 267 440 664
rect 390 255 440 267
rect 556 664 606 676
rect 556 267 562 664
rect 600 267 606 664
rect 556 255 606 267
rect -606 -267 -556 -255
rect -606 -664 -600 -267
rect -562 -664 -556 -267
rect -606 -676 -556 -664
rect -440 -267 -390 -255
rect -440 -664 -434 -267
rect -396 -664 -390 -267
rect -440 -676 -390 -664
rect -274 -267 -224 -255
rect -274 -664 -268 -267
rect -230 -664 -224 -267
rect -274 -676 -224 -664
rect -108 -267 -58 -255
rect -108 -664 -102 -267
rect -64 -664 -58 -267
rect -108 -676 -58 -664
rect 58 -267 108 -255
rect 58 -664 64 -267
rect 102 -664 108 -267
rect 58 -676 108 -664
rect 224 -267 274 -255
rect 224 -664 230 -267
rect 268 -664 274 -267
rect 224 -676 274 -664
rect 390 -267 440 -255
rect 390 -664 396 -267
rect 434 -664 440 -267
rect 390 -676 440 -664
rect 556 -267 606 -255
rect 556 -664 562 -267
rect 600 -664 606 -267
rect 556 -676 606 -664
<< res0p35 >>
rect -618 -252 -544 252
rect -452 -252 -378 252
rect -286 -252 -212 252
rect -120 -252 -46 252
rect 46 -252 120 252
rect 212 -252 286 252
rect 378 -252 452 252
rect 544 -252 618 252
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 2.5 m 1 nx 8 wmin 0.350 lmin 0.50 rho 319.8 val 3.397k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
