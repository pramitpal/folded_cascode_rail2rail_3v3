magic
tech sky130A
timestamp 1698929273
<< error_p >>
rect -54 -400 -25 400
rect 25 -400 54 400
<< mvnmos >>
rect -25 -400 25 400
<< mvndiff >>
rect -54 394 -25 400
rect -54 -394 -48 394
rect -31 -394 -25 394
rect -54 -400 -25 -394
rect 25 394 54 400
rect 25 -394 31 394
rect 48 -394 54 394
rect 25 -400 54 -394
<< mvndiffc >>
rect -48 -394 -31 394
rect 31 -394 48 394
<< poly >>
rect -25 400 25 413
rect -25 -413 25 -400
<< locali >>
rect -48 394 -31 402
rect -48 -402 -31 -394
rect 31 394 48 402
rect 31 -402 48 -394
<< viali >>
rect -48 -394 -31 394
rect 31 -394 48 394
<< metal1 >>
rect -51 394 -28 400
rect -51 -394 -48 394
rect -31 -394 -28 394
rect -51 -400 -28 -394
rect 28 394 51 400
rect 28 -394 31 394
rect 48 -394 51 394
rect 28 -400 51 -394
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
