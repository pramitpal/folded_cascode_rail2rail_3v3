magic
tech sky130A
magscale 1 2
timestamp 1697281155
<< error_p >>
rect -258 -169 -200 231
rect 200 -169 258 231
<< mvnmos >>
rect -200 -169 200 231
<< mvndiff >>
rect -258 219 -200 231
rect -258 -157 -246 219
rect -212 -157 -200 219
rect -258 -169 -200 -157
rect 200 219 258 231
rect 200 -157 212 219
rect 246 -157 258 219
rect 200 -169 258 -157
<< mvndiffc >>
rect -246 -157 -212 219
rect 212 -157 246 219
<< poly >>
rect -200 231 200 257
rect -200 -207 200 -169
rect -200 -241 -184 -207
rect 184 -241 200 -207
rect -200 -257 200 -241
<< polycont >>
rect -184 -241 184 -207
<< locali >>
rect -246 219 -212 235
rect -246 -173 -212 -157
rect 212 219 246 235
rect 212 -173 246 -157
rect -200 -241 -184 -207
rect 184 -241 200 -207
<< viali >>
rect -246 -157 -212 219
rect 212 -157 246 219
rect -184 -241 184 -207
<< metal1 >>
rect -252 219 -206 231
rect -252 -157 -246 219
rect -212 -157 -206 219
rect -252 -169 -206 -157
rect 206 219 252 231
rect 206 -157 212 219
rect 246 -157 252 219
rect 206 -169 252 -157
rect -196 -207 196 -201
rect -196 -241 -184 -207
rect 184 -241 196 -207
rect -196 -247 196 -241
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
