magic
tech sky130A
magscale 1 2
timestamp 1697284980
<< nwell >>
rect -892 -1789 1013 571
<< mvpsubdiff >>
rect -825 -2083 -777 -2036
rect -825 -3992 -818 -2083
rect -784 -3992 -777 -2083
rect 899 -2077 947 -2036
rect -825 -4020 -777 -3992
rect 899 -3986 906 -2077
rect 940 -3986 947 -2077
rect 899 -4020 947 -3986
<< mvnsubdiff >>
rect -825 352 -777 419
rect -825 -1636 -818 352
rect -784 -1636 -777 352
rect 899 390 947 419
rect -825 -1670 -777 -1636
rect 899 -1598 906 390
rect 940 -1598 947 390
rect 899 -1670 947 -1598
<< mvpsubdiffcont >>
rect -818 -3992 -784 -2083
rect 906 -3986 940 -2077
<< mvnsubdiffcont >>
rect -818 -1636 -784 352
rect 906 -1598 940 390
<< poly >>
rect -356 172 -256 219
rect -356 138 -340 172
rect -272 138 -256 172
rect -356 122 -256 138
rect -68 172 32 219
rect -68 138 -52 172
rect 16 138 32 172
rect -68 122 32 138
rect 90 172 190 219
rect 90 138 106 172
rect 174 138 190 172
rect 90 122 190 138
rect 378 172 478 219
rect 378 138 394 172
rect 462 138 478 172
rect 378 122 478 138
rect -356 -1717 -256 -1670
rect -356 -1751 -340 -1717
rect -272 -1751 -256 -1717
rect -356 -1767 -256 -1751
rect -68 -1717 32 -1670
rect -68 -1751 -52 -1717
rect 16 -1751 32 -1717
rect -68 -1767 32 -1751
rect 90 -1717 190 -1670
rect 90 -1751 106 -1717
rect 174 -1751 190 -1717
rect 90 -1767 190 -1751
rect 378 -1717 478 -1670
rect 378 -1751 394 -1717
rect 462 -1751 478 -1717
rect 378 -1767 478 -1751
rect -356 -1955 -256 -1939
rect -356 -1989 -340 -1955
rect -272 -1989 -256 -1955
rect -356 -2036 -256 -1989
rect -68 -1955 32 -1939
rect -68 -1989 -52 -1955
rect 16 -1989 32 -1955
rect -68 -2036 32 -1989
rect 90 -1955 190 -1939
rect 90 -1989 106 -1955
rect 174 -1989 190 -1955
rect 90 -2036 190 -1989
rect 378 -1955 478 -1939
rect 378 -1989 394 -1955
rect 462 -1989 478 -1955
rect 378 -2036 478 -1989
rect -356 -3848 -256 -3832
rect -356 -3882 -340 -3848
rect -272 -3882 -256 -3848
rect -356 -3920 -256 -3882
rect -68 -3848 32 -3832
rect -68 -3882 -52 -3848
rect 16 -3882 32 -3848
rect -68 -3920 32 -3882
rect 90 -3848 190 -3832
rect 90 -3882 106 -3848
rect 174 -3882 190 -3848
rect 90 -3920 190 -3882
rect 378 -3848 478 -3832
rect 378 -3882 394 -3848
rect 462 -3882 478 -3848
rect 378 -3920 478 -3882
<< polycont >>
rect -340 138 -272 172
rect -52 138 16 172
rect 106 138 174 172
rect 394 138 462 172
rect -340 -1751 -272 -1717
rect -52 -1751 16 -1717
rect 106 -1751 174 -1717
rect 394 -1751 462 -1717
rect -340 -1989 -272 -1955
rect -52 -1989 16 -1955
rect 106 -1989 174 -1955
rect 394 -1989 462 -1955
rect -340 -3882 -272 -3848
rect -52 -3882 16 -3848
rect 106 -3882 174 -3848
rect 394 -3882 462 -3848
<< locali >>
rect -690 466 812 500
rect -825 407 -777 419
rect -690 407 -656 466
rect -532 407 -498 466
rect -825 352 -656 407
rect -825 -1636 -818 352
rect -784 11 -656 352
rect -244 231 -210 466
rect 44 384 78 466
rect 332 377 366 466
rect 620 393 654 466
rect 778 407 812 466
rect 899 407 947 419
rect 778 390 947 407
rect -356 138 -340 172
rect -272 138 -52 172
rect 16 138 106 172
rect 174 138 394 172
rect 462 138 478 172
rect 44 56 599 90
rect 44 13 78 56
rect -784 -23 -498 11
rect -784 -145 -656 -23
rect -532 -87 -498 -23
rect -114 -21 236 13
rect 778 11 906 390
rect -114 -95 -80 -21
rect 202 -135 236 -21
rect 620 -23 906 11
rect 620 -138 654 -23
rect -784 -1636 -670 -145
rect -825 -1658 -670 -1636
rect 778 -1598 906 -23
rect 940 -1598 947 390
rect 982 -190 1016 56
rect 778 -1658 947 -1598
rect -825 -1670 -777 -1658
rect 899 -1670 947 -1658
rect -356 -1751 -340 -1717
rect -272 -1751 -256 -1717
rect -68 -1751 -52 -1717
rect 16 -1751 106 -1717
rect 174 -1751 190 -1717
rect 378 -1751 394 -1717
rect 462 -1751 478 -1717
rect 44 -1835 78 -1751
rect -901 -1869 78 -1835
rect 44 -1955 78 -1869
rect -356 -1989 -340 -1955
rect -272 -1989 -256 -1955
rect -68 -1989 -52 -1955
rect 16 -1989 106 -1955
rect 174 -1989 190 -1955
rect 378 -1989 394 -1955
rect 462 -1989 478 -1955
rect -825 -2048 -777 -2036
rect 899 -2048 947 -2036
rect -825 -2083 -663 -2048
rect -825 -3992 -818 -2083
rect -784 -3578 -663 -2083
rect 778 -2077 947 -2048
rect -784 -3674 -656 -3578
rect -532 -3674 -498 -3605
rect -784 -3708 -498 -3674
rect -114 -3681 -80 -3617
rect 202 -3681 236 -3604
rect -784 -3992 -656 -3708
rect -114 -3715 236 -3681
rect 620 -3674 654 -3599
rect 778 -3674 906 -2077
rect 620 -3708 906 -3674
rect 44 -3761 78 -3715
rect 44 -3795 646 -3761
rect -356 -3882 -340 -3848
rect -272 -3882 -52 -3848
rect 16 -3882 106 -3848
rect 174 -3882 394 -3848
rect 462 -3882 478 -3848
rect -825 -4008 -656 -3992
rect -825 -4020 -777 -4008
rect -690 -4058 -656 -4008
rect -532 -4058 -498 -4006
rect -244 -4058 -210 -3973
rect 44 -4058 78 -3979
rect 332 -4058 366 -3980
rect 620 -4058 654 -3959
rect 778 -3986 906 -3708
rect 940 -3986 947 -2077
rect 778 -4008 947 -3986
rect 778 -4058 812 -4008
rect 899 -4020 947 -4008
rect -690 -4092 812 -4058
<< viali >>
rect 599 56 633 90
rect 982 56 1016 90
rect -340 -1751 -272 -1717
rect 394 -1751 462 -1717
rect -340 -1989 -272 -1955
rect 394 -1989 462 -1955
rect 646 -3795 680 -3761
<< metal1 >>
rect -402 124 -368 359
rect -114 124 -80 258
rect 202 124 236 254
rect 490 124 524 254
rect -402 90 524 124
rect -401 -118 -367 90
rect -259 -30 -253 22
rect -201 -30 -195 22
rect -244 -102 -210 -30
rect 44 -119 78 90
rect 317 -30 323 22
rect 375 -30 381 22
rect 332 -111 366 -30
rect 490 -114 524 90
rect 593 90 639 102
rect 976 90 1022 102
rect 593 56 599 90
rect 633 56 982 90
rect 1016 56 1022 90
rect 593 44 639 56
rect 976 44 1022 56
rect 967 -74 973 -22
rect 1025 -74 1031 -22
rect 982 -135 1016 -74
rect -352 -1717 -260 -1711
rect 382 -1717 474 -1711
rect -352 -1751 -340 -1717
rect -272 -1751 394 -1717
rect 462 -1751 474 -1717
rect -352 -1757 -260 -1751
rect 44 -1835 78 -1751
rect 382 -1757 474 -1751
rect -874 -1869 78 -1835
rect -352 -1955 -260 -1949
rect 44 -1955 78 -1869
rect 382 -1955 474 -1949
rect -352 -1989 -340 -1955
rect -272 -1989 394 -1955
rect 462 -1989 478 -1955
rect -352 -1995 -260 -1989
rect 382 -1995 474 -1989
rect -402 -3789 -368 -3614
rect -244 -3672 -210 -3603
rect -259 -3724 -253 -3672
rect -201 -3724 -195 -3672
rect 44 -3789 78 -3601
rect 332 -3672 366 -3608
rect 317 -3724 323 -3672
rect 375 -3724 381 -3672
rect 490 -3789 524 -3589
rect -402 -3823 524 -3789
rect 640 -3761 686 -3749
rect 640 -3795 646 -3761
rect 680 -3795 1102 -3761
rect 640 -3807 686 -3795
rect -402 -3947 -368 -3823
rect -114 -3960 -80 -3823
rect 202 -3965 236 -3823
rect 490 -3945 524 -3823
<< via1 >>
rect -253 -30 -201 22
rect 323 -30 375 22
rect 973 -74 1025 -22
rect -253 -3724 -201 -3672
rect 323 -3724 375 -3672
<< metal2 >>
rect 44 56 1016 90
rect -253 22 -201 28
rect 44 13 78 56
rect 323 22 375 28
rect -201 -21 323 13
rect -253 -36 -201 -30
rect 982 -16 1016 56
rect 323 -36 375 -30
rect 973 -22 1025 -16
rect 973 -80 1025 -74
rect -253 -3672 -201 -3666
rect 323 -3672 375 -3666
rect -201 -3715 323 -3681
rect -253 -3730 -201 -3724
rect 44 -3761 78 -3715
rect 323 -3730 375 -3724
rect 44 -3795 1036 -3761
use sky130_fd_pr__nfet_g5v0d10v5_GUWUK4#0  sky130_fd_pr__nfet_g5v0d10v5_GUWUK4_0
timestamp 1697281155
transform 1 0 -594 0 1 -4001
box -108 -107 108 107
use sky130_fd_pr__nfet_g5v0d10v5_GUWUK4#0  sky130_fd_pr__nfet_g5v0d10v5_GUWUK4_1
timestamp 1697281155
transform 1 0 716 0 1 -4001
box -108 -107 108 107
use sky130_fd_pr__nfet_g5v0d10v5_SAC338  sky130_fd_pr__nfet_g5v0d10v5_SAC338_0
timestamp 1697281155
transform 1 0 -18 0 1 -2836
box -108 -826 108 826
use sky130_fd_pr__nfet_g5v0d10v5_SAC338  sky130_fd_pr__nfet_g5v0d10v5_SAC338_1
timestamp 1697281155
transform 1 0 140 0 1 -2836
box -108 -826 108 826
use sky130_fd_pr__nfet_g5v0d10v5_SAC338  sky130_fd_pr__nfet_g5v0d10v5_SAC338_2
timestamp 1697281155
transform 1 0 428 0 1 -2836
box -108 -826 108 826
use sky130_fd_pr__nfet_g5v0d10v5_SAC338  sky130_fd_pr__nfet_g5v0d10v5_SAC338_3
timestamp 1697281155
transform 1 0 -306 0 1 -2836
box -108 -826 108 826
use sky130_fd_pr__nfet_g5v0d10v5_SAT828  sky130_fd_pr__nfet_g5v0d10v5_SAT828_0
timestamp 1697281155
transform 1 0 -594 0 1 -2867
box -108 -857 108 857
use sky130_fd_pr__nfet_g5v0d10v5_SAT828  sky130_fd_pr__nfet_g5v0d10v5_SAT828_1
timestamp 1697281155
transform 1 0 716 0 1 -2867
box -108 -857 108 857
use sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0  sky130_fd_pr__nfet_g5v0d10v5_VNB5GC_0
timestamp 1697281155
transform 1 0 428 0 1 -3970
box -108 -76 108 76
use sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0  sky130_fd_pr__nfet_g5v0d10v5_VNB5GC_1
timestamp 1697281155
transform 1 0 140 0 1 -3970
box -108 -76 108 76
use sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0  sky130_fd_pr__nfet_g5v0d10v5_VNB5GC_2
timestamp 1697281155
transform 1 0 -18 0 1 -3970
box -108 -76 108 76
use sky130_fd_pr__nfet_g5v0d10v5_VNB5GC#0  sky130_fd_pr__nfet_g5v0d10v5_VNB5GC_3
timestamp 1697281155
transform 1 0 -306 0 1 -3970
box -108 -76 108 76
use sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7  sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_0
timestamp 1697284980
transform 1 0 -306 0 1 -870
box -174 -866 174 866
use sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7  sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_1
timestamp 1697284980
transform 1 0 140 0 1 -870
box -174 -866 174 866
use sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7  sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_2
timestamp 1697284980
transform 1 0 -18 0 1 -870
box -174 -866 174 866
use sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7  sky130_fd_pr__pfet_g5v0d10v5_2L5LZ7_3
timestamp 1697284980
transform 1 0 428 0 1 -870
box -174 -866 174 866
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_0
timestamp 1697281155
transform 1 0 428 0 1 319
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_1
timestamp 1697281155
transform 1 0 140 0 1 319
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_2
timestamp 1697281155
transform 1 0 -18 0 1 319
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7#0  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_3
timestamp 1697281155
transform 1 0 -306 0 1 319
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_VK4LZ7  sky130_fd_pr__pfet_g5v0d10v5_VK4LZ7_0
timestamp 1697281155
transform 1 0 -594 0 1 -834
box -174 -902 174 864
use sky130_fd_pr__pfet_g5v0d10v5_VK4LZ7  sky130_fd_pr__pfet_g5v0d10v5_VK4LZ7_1
timestamp 1697281155
transform 1 0 716 0 1 -834
box -174 -902 174 864
use sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7#0  sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_0
timestamp 1697281155
transform 1 0 -594 0 1 355
box -174 -202 174 164
use sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7#0  sky130_fd_pr__pfet_g5v0d10v5_ZUVZZ7_1
timestamp 1697281155
transform 1 0 716 0 1 355
box -174 -202 174 164
<< labels >>
flabel metal1 s -164 -1736 -164 -1736 0 FreeSans 800 0 0 0 INP
flabel locali s 59 -1815 59 -1815 0 FreeSans 800 0 0 0 INN
flabel metal2 s -164 -6 -164 -6 0 FreeSans 800 0 0 0 N3
flabel locali s 220 -37 220 -37 0 FreeSans 800 0 0 0 N4
flabel locali s -190 155 -190 155 0 FreeSans 800 0 0 0 Vb1
flabel locali s 425 483 425 483 0 FreeSans 800 0 0 0 VCC
flabel metal2 s -163 -3696 -163 -3696 0 FreeSans 800 0 0 0 N1
flabel locali s 224 -3663 224 -3663 0 FreeSans 800 0 0 0 N2
flabel locali s -149 -3863 -149 -3863 0 FreeSans 800 0 0 0 Vb5
flabel locali s 332 -4074 332 -4074 0 FreeSans 800 0 0 0 VSS
<< end >>
